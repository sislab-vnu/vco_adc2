magic
tech sky130A
timestamp 1730689382
<< locali >>
rect 245 4025 445 4035
rect 245 4005 255 4025
rect 275 4005 295 4025
rect 315 4005 335 4025
rect 355 4005 375 4025
rect 395 4005 415 4025
rect 435 4005 445 4025
rect 245 3995 445 4005
rect 2110 4025 2310 4035
rect 2110 4005 2120 4025
rect 2140 4005 2160 4025
rect 2180 4005 2200 4025
rect 2220 4005 2240 4025
rect 2260 4005 2280 4025
rect 2300 4005 2310 4025
rect 2110 3995 2310 4005
rect 565 -780 3055 -770
rect 565 -800 575 -780
rect 595 -800 615 -780
rect 635 -800 2985 -780
rect 3005 -800 3025 -780
rect 3045 -800 3055 -780
rect 565 -810 3055 -800
rect 3015 -820 3055 -810
rect 3015 -840 3025 -820
rect 3045 -840 3055 -820
rect 3015 -850 3055 -840
rect 735 -1075 1370 -1065
rect 735 -1105 1210 -1075
rect 1240 -1105 1270 -1075
rect 1300 -1105 1330 -1075
rect 1360 -1105 1370 -1075
rect 735 -1110 1370 -1105
rect 765 -1115 1370 -1110
rect -1120 -3375 -915 -3370
rect -1120 -3380 -910 -3375
rect -1120 -3400 -1110 -3380
rect -1090 -3400 -1070 -3380
rect -1050 -3400 -910 -3380
rect -1120 -3410 -910 -3400
rect -1120 -3420 -1080 -3410
rect -1120 -3440 -1110 -3420
rect -1090 -3440 -1080 -3420
rect -1120 -3450 -1080 -3440
rect 630 -3945 1185 -3935
rect 630 -3965 640 -3945
rect 660 -3965 680 -3945
rect 700 -3965 720 -3945
rect 740 -3965 1075 -3945
rect 1095 -3965 1115 -3945
rect 1135 -3965 1155 -3945
rect 1175 -3965 1185 -3945
rect 630 -3975 1185 -3965
rect 8140 -3950 8585 -3935
rect 8140 -3970 8155 -3950
rect 8175 -3970 8195 -3950
rect 8215 -3970 8585 -3950
rect 8140 -3985 8585 -3970
rect 8140 -3990 8190 -3985
rect 8140 -4010 8155 -3990
rect 8175 -4010 8190 -3990
rect 8140 -4025 8190 -4010
rect -820 -4570 -690 -4550
rect -1420 -4590 -690 -4570
rect -1420 -4620 -1400 -4590
rect -1370 -4620 -1340 -4590
rect -1310 -4620 -690 -4590
rect -1420 -4650 -690 -4620
rect -1420 -4680 -1400 -4650
rect -1370 -4680 -1340 -4650
rect -1310 -4680 -690 -4650
rect -1420 -4690 -690 -4680
rect 8535 -4980 8585 -3985
rect 8535 -5000 8550 -4980
rect 8570 -5000 8585 -4980
rect 8535 -5010 8585 -5000
rect 8500 -5020 8585 -5010
rect 8500 -5040 8510 -5020
rect 8530 -5040 8550 -5020
rect 8570 -5040 8585 -5020
rect 8500 -5050 8585 -5040
<< viali >>
rect 255 4005 275 4025
rect 295 4005 315 4025
rect 335 4005 355 4025
rect 375 4005 395 4025
rect 415 4005 435 4025
rect 2120 4005 2140 4025
rect 2160 4005 2180 4025
rect 2200 4005 2220 4025
rect 2240 4005 2260 4025
rect 2280 4005 2300 4025
rect 5530 4005 5550 4025
rect 5570 4005 5590 4025
rect 5610 4005 5630 4025
rect 5650 4005 5670 4025
rect 5690 4005 5710 4025
rect 7945 4005 7965 4025
rect 7985 4005 8005 4025
rect 8025 4005 8045 4025
rect 8065 4005 8085 4025
rect 8105 4005 8125 4025
rect -1000 -235 -980 -215
rect -960 -235 -940 -215
rect 575 -800 595 -780
rect 615 -800 635 -780
rect 2985 -800 3005 -780
rect 3025 -800 3045 -780
rect 3025 -840 3045 -820
rect 1210 -1105 1240 -1075
rect 1270 -1105 1300 -1075
rect 1330 -1105 1360 -1075
rect -1110 -3400 -1090 -3380
rect -1070 -3400 -1050 -3380
rect -1110 -3440 -1090 -3420
rect 640 -3965 660 -3945
rect 680 -3965 700 -3945
rect 720 -3965 740 -3945
rect 1075 -3965 1095 -3945
rect 1115 -3965 1135 -3945
rect 1155 -3965 1175 -3945
rect 8155 -3970 8175 -3950
rect 8195 -3970 8215 -3950
rect 8155 -4010 8175 -3990
rect -1400 -4620 -1370 -4590
rect -1340 -4620 -1310 -4590
rect -1400 -4680 -1370 -4650
rect -1340 -4680 -1310 -4650
rect 8550 -5000 8570 -4980
rect 8510 -5040 8530 -5020
rect 8550 -5040 8570 -5020
<< metal1 >>
rect 245 4030 445 4035
rect 245 4000 250 4030
rect 280 4025 310 4030
rect 340 4025 370 4030
rect 400 4025 445 4030
rect 280 4005 295 4025
rect 355 4005 370 4025
rect 400 4005 415 4025
rect 435 4005 445 4025
rect 280 4000 310 4005
rect 340 4000 370 4005
rect 400 4000 445 4005
rect 245 3995 445 4000
rect 2110 4030 2310 4035
rect 2110 4000 2115 4030
rect 2145 4025 2195 4030
rect 2225 4025 2275 4030
rect 2145 4005 2160 4025
rect 2180 4005 2195 4025
rect 2225 4005 2240 4025
rect 2260 4005 2275 4025
rect 2145 4000 2195 4005
rect 2225 4000 2275 4005
rect 2305 4000 2310 4030
rect 2110 3995 2310 4000
rect 5520 4030 5720 4035
rect 5520 4000 5525 4030
rect 5555 4025 5605 4030
rect 5635 4025 5685 4030
rect 5555 4005 5570 4025
rect 5590 4005 5605 4025
rect 5635 4005 5650 4025
rect 5670 4005 5685 4025
rect 5555 4000 5605 4005
rect 5635 4000 5685 4005
rect 5715 4000 5720 4030
rect 5520 3995 5720 4000
rect 7935 4030 8135 4035
rect 7935 4000 7940 4030
rect 7970 4025 8020 4030
rect 8050 4025 8100 4030
rect 7970 4005 7985 4025
rect 8005 4005 8020 4025
rect 8050 4005 8065 4025
rect 8085 4005 8100 4025
rect 7970 4000 8020 4005
rect 8050 4000 8100 4005
rect 8130 4000 8135 4030
rect 7935 3995 8135 4000
rect 3445 2450 3570 2480
rect 3445 2420 3455 2450
rect 3485 2420 3515 2450
rect 3545 2420 3570 2450
rect 3445 2400 3570 2420
rect -1010 -205 -960 1050
rect -740 540 -540 555
rect -740 505 -715 540
rect -680 505 -600 540
rect -565 505 -540 540
rect -740 -65 -540 505
rect -160 535 40 555
rect -160 500 -135 535
rect -100 500 -25 535
rect 10 500 40 535
rect -160 -60 40 500
rect 445 540 645 555
rect 445 510 465 540
rect 495 510 590 540
rect 620 510 645 540
rect 445 -65 645 510
rect -1010 -215 -930 -205
rect -1010 -235 -1000 -215
rect -980 -235 -960 -215
rect -940 -235 -930 -215
rect -1010 -245 -930 -235
rect 485 -780 645 -770
rect 485 -800 575 -780
rect 595 -800 615 -780
rect 635 -800 645 -780
rect 485 -810 645 -800
rect 2975 -780 3055 -770
rect 2975 -800 2985 -780
rect 3005 -800 3025 -780
rect 3045 -800 3055 -780
rect 2975 -810 3055 -800
rect 3015 -820 3055 -810
rect 3015 -840 3025 -820
rect 3045 -840 3055 -820
rect 1200 -1075 1370 -1065
rect 1200 -1105 1210 -1075
rect 1240 -1105 1270 -1075
rect 1300 -1105 1330 -1075
rect 1360 -1105 1370 -1075
rect 1200 -1115 1370 -1105
rect 1180 -1550 1380 -1115
rect 1180 -1580 1195 -1550
rect 1225 -1580 1255 -1550
rect 1285 -1580 1315 -1550
rect 1345 -1580 1380 -1550
rect 1180 -1610 1380 -1580
rect 1180 -1640 1195 -1610
rect 1225 -1640 1255 -1610
rect 1285 -1640 1315 -1610
rect 1345 -1640 1380 -1610
rect 1180 -1740 1380 -1640
rect -1160 -2245 -960 -1950
rect -1160 -2275 -1140 -2245
rect -1110 -2275 -1015 -2245
rect -985 -2275 -960 -2245
rect -1160 -2400 -960 -2275
rect 3015 -2415 3055 -840
rect 9255 -1205 9305 -1170
rect 9255 -1235 9265 -1205
rect 9295 -1235 9305 -1205
rect 9255 -1265 9305 -1235
rect 9255 -1295 9265 -1265
rect 9295 -1295 9305 -1265
rect 9255 -1325 9305 -1295
rect 9255 -1355 9265 -1325
rect 9295 -1355 9305 -1325
rect 9255 -1370 9305 -1355
rect 6580 -1790 6625 -1770
rect 6580 -1820 6585 -1790
rect 6615 -1820 6625 -1790
rect 6580 -1850 6625 -1820
rect 6580 -1880 6585 -1850
rect 6615 -1880 6625 -1850
rect 6580 -1945 6625 -1880
rect 3500 -2210 3610 -2200
rect 3500 -2240 3510 -2210
rect 3540 -2240 3570 -2210
rect 3600 -2240 3610 -2210
rect 3500 -2250 3610 -2240
rect 3500 -2270 4120 -2250
rect 3500 -2300 3510 -2270
rect 3540 -2300 3570 -2270
rect 3600 -2300 4120 -2270
rect 3500 -2310 3610 -2300
rect 3015 -2455 3260 -2415
rect -895 -3035 -855 -2510
rect -740 -2750 -540 -2670
rect -740 -2780 -725 -2750
rect -695 -2780 -665 -2750
rect -635 -2780 -605 -2750
rect -575 -2780 -540 -2750
rect -740 -2790 -540 -2780
rect 125 -2750 325 -2665
rect 125 -2780 140 -2750
rect 170 -2780 200 -2750
rect 230 -2780 260 -2750
rect 290 -2780 325 -2750
rect 125 -2790 325 -2780
rect 1045 -2750 1245 -2665
rect 1045 -2780 1060 -2750
rect 1090 -2780 1120 -2750
rect 1150 -2780 1180 -2750
rect 1210 -2780 1245 -2750
rect 1045 -2790 1245 -2780
rect -895 -3075 1185 -3035
rect -1120 -3380 -1040 -3370
rect -1120 -3400 -1110 -3380
rect -1090 -3400 -1070 -3380
rect -1050 -3400 -1040 -3380
rect -1120 -3410 -1040 -3400
rect -1120 -3420 -1080 -3410
rect -1120 -3440 -1110 -3420
rect -1090 -3440 -1080 -3420
rect -1620 -4585 -1300 -4570
rect -1620 -4615 -1605 -4585
rect -1575 -4615 -1545 -4585
rect -1515 -4615 -1485 -4585
rect -1455 -4590 -1300 -4585
rect -1455 -4615 -1400 -4590
rect -1620 -4620 -1400 -4615
rect -1370 -4620 -1340 -4590
rect -1310 -4620 -1300 -4590
rect -1620 -4650 -1300 -4620
rect -1620 -4680 -1400 -4650
rect -1370 -4680 -1340 -4650
rect -1310 -4680 -1300 -4650
rect -1620 -4685 -1300 -4680
rect -1420 -4690 -1300 -4685
rect -1120 -5010 -1080 -3440
rect -980 -3545 -740 -3530
rect -980 -3575 -965 -3545
rect -935 -3575 -905 -3545
rect -875 -3575 -845 -3545
rect -815 -3575 -785 -3545
rect -755 -3575 -740 -3545
rect -980 -3585 -740 -3575
rect 1145 -3935 1185 -3075
rect 3220 -3505 3260 -2455
rect 4555 -2475 4655 -2465
rect 4555 -2505 4565 -2475
rect 4595 -2505 4615 -2475
rect 4645 -2505 4655 -2475
rect 4555 -2525 4655 -2505
rect 4555 -2555 4565 -2525
rect 4595 -2555 4615 -2525
rect 4645 -2555 4655 -2525
rect 4555 -2565 4655 -2555
rect 485 -3945 750 -3935
rect 485 -3965 640 -3945
rect 660 -3965 680 -3945
rect 700 -3965 720 -3945
rect 740 -3965 750 -3945
rect 485 -3975 750 -3965
rect 1065 -3945 1185 -3935
rect 1065 -3965 1075 -3945
rect 1095 -3965 1115 -3945
rect 1135 -3965 1155 -3945
rect 1175 -3965 1185 -3945
rect 1065 -3975 1185 -3965
rect 8140 -3950 8245 -3935
rect 8140 -3970 8155 -3950
rect 8175 -3970 8195 -3950
rect 8215 -3970 8245 -3950
rect 8140 -3985 8245 -3970
rect 8140 -3990 8190 -3985
rect 8140 -4010 8155 -3990
rect 8175 -4010 8190 -3990
rect 8140 -4025 8190 -4010
rect 6125 -4070 6325 -4060
rect 6125 -4100 6140 -4070
rect 6170 -4100 6200 -4070
rect 6230 -4100 6260 -4070
rect 6290 -4100 6325 -4070
rect 6125 -4110 6325 -4100
rect -820 -4570 -620 -4525
rect 290 -4580 490 -4530
rect 290 -4610 305 -4580
rect 335 -4610 365 -4580
rect 395 -4610 425 -4580
rect 455 -4610 490 -4580
rect 290 -4625 490 -4610
rect 8535 -4980 8585 -4970
rect 8535 -5000 8550 -4980
rect 8570 -5000 8585 -4980
rect 8535 -5010 8585 -5000
rect -1120 -5020 8585 -5010
rect -1120 -5040 8510 -5020
rect 8530 -5040 8550 -5020
rect 8570 -5040 8585 -5020
rect -1120 -5050 8585 -5040
<< via1 >>
rect 250 4025 280 4030
rect 310 4025 340 4030
rect 370 4025 400 4030
rect 250 4005 255 4025
rect 255 4005 275 4025
rect 275 4005 280 4025
rect 310 4005 315 4025
rect 315 4005 335 4025
rect 335 4005 340 4025
rect 370 4005 375 4025
rect 375 4005 395 4025
rect 395 4005 400 4025
rect 250 4000 280 4005
rect 310 4000 340 4005
rect 370 4000 400 4005
rect 2115 4025 2145 4030
rect 2195 4025 2225 4030
rect 2275 4025 2305 4030
rect 2115 4005 2120 4025
rect 2120 4005 2140 4025
rect 2140 4005 2145 4025
rect 2195 4005 2200 4025
rect 2200 4005 2220 4025
rect 2220 4005 2225 4025
rect 2275 4005 2280 4025
rect 2280 4005 2300 4025
rect 2300 4005 2305 4025
rect 2115 4000 2145 4005
rect 2195 4000 2225 4005
rect 2275 4000 2305 4005
rect 5525 4025 5555 4030
rect 5605 4025 5635 4030
rect 5685 4025 5715 4030
rect 5525 4005 5530 4025
rect 5530 4005 5550 4025
rect 5550 4005 5555 4025
rect 5605 4005 5610 4025
rect 5610 4005 5630 4025
rect 5630 4005 5635 4025
rect 5685 4005 5690 4025
rect 5690 4005 5710 4025
rect 5710 4005 5715 4025
rect 5525 4000 5555 4005
rect 5605 4000 5635 4005
rect 5685 4000 5715 4005
rect 7940 4025 7970 4030
rect 8020 4025 8050 4030
rect 8100 4025 8130 4030
rect 7940 4005 7945 4025
rect 7945 4005 7965 4025
rect 7965 4005 7970 4025
rect 8020 4005 8025 4025
rect 8025 4005 8045 4025
rect 8045 4005 8050 4025
rect 8100 4005 8105 4025
rect 8105 4005 8125 4025
rect 8125 4005 8130 4025
rect 7940 4000 7970 4005
rect 8020 4000 8050 4005
rect 8100 4000 8130 4005
rect 3455 2420 3485 2450
rect 3515 2420 3545 2450
rect 7350 2285 7380 2315
rect 7350 2225 7380 2255
rect 7350 2165 7380 2195
rect -715 505 -680 540
rect -600 505 -565 540
rect -135 500 -100 535
rect -25 500 10 535
rect 465 510 495 540
rect 590 510 620 540
rect 1195 -1580 1225 -1550
rect 1255 -1580 1285 -1550
rect 1315 -1580 1345 -1550
rect 1195 -1640 1225 -1610
rect 1255 -1640 1285 -1610
rect 1315 -1640 1345 -1610
rect -1140 -2275 -1110 -2245
rect -1015 -2275 -985 -2245
rect 9265 -1235 9295 -1205
rect 9265 -1295 9295 -1265
rect 9265 -1355 9295 -1325
rect 6585 -1820 6615 -1790
rect 6585 -1880 6615 -1850
rect 3510 -2240 3540 -2210
rect 3570 -2240 3600 -2210
rect 3510 -2300 3540 -2270
rect 3570 -2300 3600 -2270
rect -725 -2780 -695 -2750
rect -665 -2780 -635 -2750
rect -605 -2780 -575 -2750
rect 140 -2780 170 -2750
rect 200 -2780 230 -2750
rect 260 -2780 290 -2750
rect 1060 -2780 1090 -2750
rect 1120 -2780 1150 -2750
rect 1180 -2780 1210 -2750
rect -1605 -4615 -1575 -4585
rect -1545 -4615 -1515 -4585
rect -1485 -4615 -1455 -4585
rect -965 -3575 -935 -3545
rect -905 -3575 -875 -3545
rect -845 -3575 -815 -3545
rect -785 -3575 -755 -3545
rect 4565 -2505 4595 -2475
rect 4615 -2505 4645 -2475
rect 4565 -2555 4595 -2525
rect 4615 -2555 4645 -2525
rect 9265 -3535 9295 -3505
rect 9265 -3595 9295 -3565
rect 9265 -3655 9295 -3625
rect 6140 -4100 6170 -4070
rect 6200 -4100 6230 -4070
rect 6260 -4100 6290 -4070
rect 305 -4610 335 -4580
rect 365 -4610 395 -4580
rect 425 -4610 455 -4580
rect 4015 -4820 4045 -4790
rect 4075 -4820 4105 -4790
rect 4135 -4820 4165 -4790
rect 8045 -4820 8075 -4790
rect 8105 -4820 8135 -4790
rect 8165 -4820 8195 -4790
<< metal2 >>
rect 21030 16365 21370 16765
rect 20245 16165 21370 16365
rect -7675 12995 -3415 13035
rect -7675 12895 -7615 12995
rect -7515 12895 -7415 12995
rect -7315 12895 -7215 12995
rect -7115 12895 -3415 12995
rect -7675 12835 -3415 12895
rect -3615 -1810 -3415 12835
rect 245 4090 445 4105
rect 245 4050 265 4090
rect 305 4050 385 4090
rect 425 4050 445 4090
rect 245 4030 445 4050
rect 245 4000 250 4030
rect 280 4000 310 4030
rect 340 4000 370 4030
rect 400 4000 445 4030
rect 245 3995 445 4000
rect 2110 4095 2310 4105
rect 2110 4055 2130 4095
rect 2170 4055 2240 4095
rect 2280 4055 2310 4095
rect 2110 4030 2310 4055
rect 2110 4000 2115 4030
rect 2145 4000 2195 4030
rect 2225 4000 2275 4030
rect 2305 4000 2310 4030
rect 2110 3995 2310 4000
rect 5520 4095 5720 4110
rect 5520 4055 5540 4095
rect 5580 4055 5655 4095
rect 5695 4055 5720 4095
rect 5520 4030 5720 4055
rect 5520 4000 5525 4030
rect 5555 4000 5605 4030
rect 5635 4000 5685 4030
rect 5715 4000 5720 4030
rect 5520 3995 5720 4000
rect 7935 4090 8135 4105
rect 7935 4050 7950 4090
rect 7990 4050 8070 4090
rect 8110 4050 8135 4090
rect 7935 4030 8135 4050
rect 7935 4000 7940 4030
rect 7970 4000 8020 4030
rect 8050 4000 8100 4030
rect 8130 4000 8135 4030
rect 7935 3995 8135 4000
rect 20245 2550 20445 16165
rect 21030 15835 21370 16165
rect 11245 2500 20445 2550
rect 3570 2480 20445 2500
rect 3445 2450 20445 2480
rect 3445 2420 3455 2450
rect 3485 2420 3515 2450
rect 3545 2420 20445 2450
rect 3445 2400 20445 2420
rect 11245 2350 20445 2400
rect 7340 2320 7495 2350
rect 7340 2315 7415 2320
rect 7340 2285 7350 2315
rect 7380 2285 7415 2315
rect 7340 2270 7415 2285
rect 7465 2270 7495 2320
rect 7340 2255 7495 2270
rect 7340 2225 7350 2255
rect 7380 2225 7495 2255
rect 7340 2220 7495 2225
rect 7340 2195 7415 2220
rect 7340 2165 7350 2195
rect 7380 2170 7415 2195
rect 7465 2170 7495 2220
rect 7380 2165 7495 2170
rect 7340 2150 7495 2165
rect -740 540 -540 555
rect -740 505 -715 540
rect -680 505 -600 540
rect -565 505 -540 540
rect -740 480 -540 505
rect -740 440 -715 480
rect -675 440 -610 480
rect -570 440 -540 480
rect -740 410 -540 440
rect -740 370 -715 410
rect -675 370 -610 410
rect -570 370 -540 410
rect -740 355 -540 370
rect -160 535 40 555
rect -160 500 -135 535
rect -100 500 -25 535
rect 10 500 40 535
rect -160 475 40 500
rect -160 435 -135 475
rect -95 435 -25 475
rect 15 435 40 475
rect -160 405 40 435
rect -160 365 -135 405
rect -95 365 -25 405
rect 15 365 40 405
rect -160 355 40 365
rect 445 540 645 555
rect 445 510 465 540
rect 495 510 590 540
rect 620 510 645 540
rect 445 490 645 510
rect 445 450 465 490
rect 505 450 585 490
rect 625 450 645 490
rect 445 410 645 450
rect 445 370 465 410
rect 505 370 585 410
rect 625 370 645 410
rect 445 355 645 370
rect 9255 -1195 9395 -1170
rect 9255 -1205 9325 -1195
rect 9255 -1235 9265 -1205
rect 9295 -1235 9325 -1205
rect 9365 -1235 9395 -1195
rect 9255 -1265 9395 -1235
rect 9255 -1295 9265 -1265
rect 9295 -1275 9395 -1265
rect 9295 -1295 9325 -1275
rect 9255 -1315 9325 -1295
rect 9365 -1315 9395 -1275
rect 9255 -1325 9395 -1315
rect 9255 -1355 9265 -1325
rect 9295 -1355 9395 -1325
rect 9255 -1370 9395 -1355
rect 1180 -1550 1380 -1540
rect 1180 -1580 1195 -1550
rect 1225 -1580 1255 -1550
rect 1285 -1580 1315 -1550
rect 1345 -1580 1380 -1550
rect 1180 -1610 1380 -1580
rect 1180 -1640 1195 -1610
rect 1225 -1640 1255 -1610
rect 1285 -1640 1315 -1610
rect 1345 -1640 1380 -1610
rect 1180 -1670 1380 -1640
rect 1180 -1710 1190 -1670
rect 1230 -1710 1270 -1670
rect 1310 -1710 1380 -1670
rect 1180 -1715 1380 -1710
rect 6580 -1785 6710 -1770
rect 6580 -1790 6650 -1785
rect -3615 -1920 2510 -1810
rect -1160 -2110 -960 -2095
rect -1160 -2150 -1145 -2110
rect -1105 -2150 -1020 -2110
rect -980 -2150 -960 -2110
rect -1160 -2185 -960 -2150
rect -1160 -2225 -1145 -2185
rect -1105 -2225 -1020 -2185
rect -980 -2225 -960 -2185
rect -1160 -2245 -960 -2225
rect -1160 -2275 -1140 -2245
rect -1110 -2275 -1015 -2245
rect -985 -2275 -960 -2245
rect -1160 -2295 -960 -2275
rect 2400 -2200 2510 -1920
rect 6580 -1820 6585 -1790
rect 6615 -1820 6650 -1790
rect 6580 -1825 6650 -1820
rect 6690 -1825 6710 -1785
rect 6580 -1850 6710 -1825
rect 6580 -1880 6585 -1850
rect 6615 -1880 6710 -1850
rect 6580 -1905 6710 -1880
rect 6580 -1945 6650 -1905
rect 6690 -1945 6710 -1905
rect 6580 -1970 6710 -1945
rect 2400 -2210 3610 -2200
rect 2400 -2240 3510 -2210
rect 3540 -2240 3570 -2210
rect 3600 -2240 3610 -2210
rect 2400 -2270 3610 -2240
rect 2400 -2300 3510 -2270
rect 3540 -2300 3570 -2270
rect 3600 -2300 3610 -2270
rect 2400 -2310 3610 -2300
rect 4555 -2475 4655 -2465
rect 4555 -2505 4565 -2475
rect 4595 -2505 4615 -2475
rect 4645 -2505 4655 -2475
rect 4555 -2525 4655 -2505
rect 4555 -2555 4565 -2525
rect 4595 -2555 4615 -2525
rect 4645 -2555 4655 -2525
rect -740 -2750 -540 -2735
rect -740 -2780 -725 -2750
rect -695 -2780 -665 -2750
rect -635 -2780 -605 -2750
rect -575 -2780 -540 -2750
rect -740 -2815 -540 -2780
rect -740 -2855 -715 -2815
rect -675 -2855 -615 -2815
rect -575 -2855 -540 -2815
rect -740 -2885 -540 -2855
rect -740 -2925 -715 -2885
rect -675 -2925 -615 -2885
rect -575 -2925 -540 -2885
rect -740 -2935 -540 -2925
rect 125 -2750 325 -2735
rect 125 -2780 140 -2750
rect 170 -2780 200 -2750
rect 230 -2780 260 -2750
rect 290 -2780 325 -2750
rect 125 -2815 325 -2780
rect 125 -2855 150 -2815
rect 190 -2855 250 -2815
rect 290 -2855 325 -2815
rect 125 -2885 325 -2855
rect 125 -2925 150 -2885
rect 190 -2925 250 -2885
rect 290 -2925 325 -2885
rect 125 -2935 325 -2925
rect 1045 -2750 1245 -2735
rect 1045 -2780 1060 -2750
rect 1090 -2780 1120 -2750
rect 1150 -2780 1180 -2750
rect 1210 -2780 1245 -2750
rect 1045 -2815 1245 -2780
rect 1045 -2855 1070 -2815
rect 1110 -2855 1170 -2815
rect 1210 -2855 1245 -2815
rect 1045 -2885 1245 -2855
rect 4555 -2860 4655 -2555
rect 1045 -2925 1070 -2885
rect 1110 -2925 1170 -2885
rect 1210 -2925 1245 -2885
rect 1045 -2935 1245 -2925
rect 3530 -2960 4655 -2860
rect -980 -3545 -740 -3530
rect -980 -3575 -965 -3545
rect -935 -3575 -905 -3545
rect -875 -3575 -845 -3545
rect -815 -3575 -785 -3545
rect -755 -3575 -740 -3545
rect -980 -3605 -740 -3575
rect -980 -3645 -965 -3605
rect -925 -3645 -885 -3605
rect -845 -3645 -805 -3605
rect -765 -3645 -740 -3605
rect -980 -3660 -740 -3645
rect -1620 -4585 -1420 -4575
rect -1620 -4615 -1605 -4585
rect -1575 -4615 -1545 -4585
rect -1515 -4615 -1485 -4585
rect -1455 -4615 -1420 -4585
rect -1620 -4630 -1420 -4615
rect -1620 -4670 -1605 -4630
rect -1565 -4670 -1490 -4630
rect -1450 -4670 -1420 -4630
rect -1620 -4685 -1420 -4670
rect 290 -4580 490 -4570
rect 290 -4610 305 -4580
rect 335 -4610 365 -4580
rect 395 -4610 425 -4580
rect 455 -4610 490 -4580
rect 290 -4630 490 -4610
rect 290 -4670 305 -4630
rect 345 -4670 420 -4630
rect 460 -4670 490 -4630
rect 290 -4680 490 -4670
rect 3530 -8600 3730 -2960
rect 9255 -3505 9380 -3470
rect 9255 -3535 9265 -3505
rect 9295 -3535 9380 -3505
rect 9255 -3565 9325 -3535
rect 9255 -3595 9265 -3565
rect 9295 -3575 9325 -3565
rect 9365 -3575 9380 -3535
rect 9295 -3595 9380 -3575
rect 9255 -3615 9380 -3595
rect 9255 -3625 9325 -3615
rect 9255 -3655 9265 -3625
rect 9295 -3655 9325 -3625
rect 9365 -3655 9380 -3615
rect 9255 -3670 9380 -3655
rect 6125 -4070 6325 -4060
rect 6125 -4100 6140 -4070
rect 6170 -4100 6200 -4070
rect 6230 -4100 6260 -4070
rect 6290 -4100 6325 -4070
rect 6125 -4115 6325 -4100
rect 6125 -4155 6135 -4115
rect 6175 -4155 6255 -4115
rect 6295 -4155 6325 -4115
rect 6125 -4160 6325 -4155
rect 4000 -4790 4195 -4780
rect 4000 -4820 4015 -4790
rect 4045 -4820 4075 -4790
rect 4105 -4820 4135 -4790
rect 4165 -4820 4195 -4790
rect 4000 -4845 4195 -4820
rect 4000 -4885 4020 -4845
rect 4060 -4885 4130 -4845
rect 4170 -4885 4195 -4845
rect 4000 -4900 4195 -4885
rect 8035 -4790 8230 -4780
rect 8035 -4820 8045 -4790
rect 8075 -4820 8105 -4790
rect 8135 -4820 8165 -4790
rect 8195 -4820 8230 -4790
rect 8035 -4845 8230 -4820
rect 8035 -4885 8050 -4845
rect 8090 -4885 8170 -4845
rect 8210 -4885 8230 -4845
rect 8035 -4900 8230 -4885
rect -5410 -8800 3730 -8600
rect -5410 -13085 -5210 -9130
rect -7645 -13150 -5210 -13085
rect -7645 -13220 -7595 -13150
rect -7525 -13220 -7455 -13150
rect -7385 -13220 -7315 -13150
rect -7245 -13220 -7175 -13150
rect -7105 -13220 -7040 -13150
rect -6970 -13220 -5210 -13150
rect -7645 -13285 -5210 -13220
<< via2 >>
rect -7615 12895 -7515 12995
rect -7415 12895 -7315 12995
rect -7215 12895 -7115 12995
rect 265 4050 305 4090
rect 385 4050 425 4090
rect 2130 4055 2170 4095
rect 2240 4055 2280 4095
rect 5540 4055 5580 4095
rect 5655 4055 5695 4095
rect 7950 4050 7990 4090
rect 8070 4050 8110 4090
rect 7415 2270 7465 2320
rect 7415 2170 7465 2220
rect -715 440 -675 480
rect -610 440 -570 480
rect -715 370 -675 410
rect -610 370 -570 410
rect -135 435 -95 475
rect -25 435 15 475
rect -135 365 -95 405
rect -25 365 15 405
rect 465 450 505 490
rect 585 450 625 490
rect 465 370 505 410
rect 585 370 625 410
rect 9325 -1235 9365 -1195
rect 9325 -1315 9365 -1275
rect 1190 -1710 1230 -1670
rect 1270 -1710 1310 -1670
rect -1145 -2150 -1105 -2110
rect -1020 -2150 -980 -2110
rect -1145 -2225 -1105 -2185
rect -1020 -2225 -980 -2185
rect 6650 -1825 6690 -1785
rect 6650 -1945 6690 -1905
rect -715 -2855 -675 -2815
rect -615 -2855 -575 -2815
rect -715 -2925 -675 -2885
rect -615 -2925 -575 -2885
rect 150 -2855 190 -2815
rect 250 -2855 290 -2815
rect 150 -2925 190 -2885
rect 250 -2925 290 -2885
rect 1070 -2855 1110 -2815
rect 1170 -2855 1210 -2815
rect 1070 -2925 1110 -2885
rect 1170 -2925 1210 -2885
rect -965 -3645 -925 -3605
rect -885 -3645 -845 -3605
rect -805 -3645 -765 -3605
rect -1605 -4670 -1565 -4630
rect -1490 -4670 -1450 -4630
rect 305 -4670 345 -4630
rect 420 -4670 460 -4630
rect 9325 -3575 9365 -3535
rect 9325 -3655 9365 -3615
rect 6135 -4155 6175 -4115
rect 6255 -4155 6295 -4115
rect 4020 -4885 4060 -4845
rect 4130 -4885 4170 -4845
rect 8050 -4885 8090 -4845
rect 8170 -4885 8210 -4845
rect -7595 -13220 -7525 -13150
rect -7455 -13220 -7385 -13150
rect -7315 -13220 -7245 -13150
rect -7175 -13220 -7105 -13150
rect -7040 -13220 -6970 -13150
<< metal3 >>
rect -7675 12995 -6965 13035
rect -7675 12895 -7615 12995
rect -7515 12895 -7415 12995
rect -7315 12895 -7215 12995
rect -7115 12895 -6965 12995
rect -7675 12835 -6965 12895
rect -3162 5905 11050 5950
rect -3162 5870 265 5905
rect -3162 5820 -3120 5870
rect -3070 5820 -3020 5870
rect -2970 5855 265 5870
rect 315 5855 365 5905
rect 415 5890 11050 5905
rect 415 5855 2130 5890
rect -2970 5840 2130 5855
rect 2180 5840 2230 5890
rect 2280 5870 11050 5890
rect 2280 5865 7960 5870
rect 2280 5840 5540 5865
rect -2970 5820 5540 5840
rect -3162 5815 5540 5820
rect 5590 5815 5640 5865
rect 5690 5820 7960 5865
rect 8010 5820 8060 5870
rect 8110 5865 11050 5870
rect 8110 5820 10810 5865
rect 5690 5815 10810 5820
rect 10860 5815 10910 5865
rect 10960 5815 11050 5865
rect -3162 5805 11050 5815
rect -3162 5770 265 5805
rect -3162 5720 -3120 5770
rect -3070 5720 -3020 5770
rect -2970 5755 265 5770
rect 315 5755 365 5805
rect 415 5790 11050 5805
rect 415 5755 2130 5790
rect -2970 5740 2130 5755
rect 2180 5740 2230 5790
rect 2280 5770 11050 5790
rect 2280 5765 7960 5770
rect 2280 5740 5540 5765
rect -2970 5720 5540 5740
rect -3162 5715 5540 5720
rect 5590 5715 5640 5765
rect 5690 5720 7960 5765
rect 8010 5720 8060 5770
rect 8110 5765 11050 5770
rect 8110 5720 10810 5765
rect 5690 5715 10810 5720
rect 10860 5715 10910 5765
rect 10960 5715 11050 5765
rect -3162 5678 11050 5715
rect -565 5675 -340 5678
rect -2074 4870 10030 4930
rect -2074 4820 -2035 4870
rect -1985 4820 -1935 4870
rect -1885 4865 10030 4870
rect -1885 4820 9850 4865
rect -2074 4815 9850 4820
rect 9900 4815 9950 4865
rect 10000 4815 10030 4865
rect -2074 4770 10030 4815
rect -2074 4720 -2035 4770
rect -1985 4720 -1935 4770
rect -1885 4765 10030 4770
rect -1885 4720 9850 4765
rect -2074 4715 9850 4720
rect 9900 4715 9950 4765
rect 10000 4715 10030 4765
rect -2074 4658 10030 4715
rect 245 4175 445 4185
rect 245 4125 265 4175
rect 315 4125 365 4175
rect 415 4125 445 4175
rect 245 4100 445 4125
rect 245 4040 255 4100
rect 315 4040 375 4100
rect 435 4040 445 4100
rect 245 4035 445 4040
rect 2110 4175 2310 4185
rect 2110 4125 2130 4175
rect 2180 4125 2230 4175
rect 2280 4125 2310 4175
rect 2110 4095 2310 4125
rect 2110 4055 2130 4095
rect 2170 4055 2240 4095
rect 2280 4055 2310 4095
rect 2110 4035 2310 4055
rect 5520 4175 5720 4185
rect 5520 4125 5540 4175
rect 5590 4125 5640 4175
rect 5690 4125 5720 4175
rect 5520 4095 5720 4125
rect 5520 4055 5540 4095
rect 5580 4055 5655 4095
rect 5695 4055 5720 4095
rect 5520 4035 5720 4055
rect 7935 4165 8135 4175
rect 7935 4115 7950 4165
rect 8000 4115 8065 4165
rect 8115 4115 8135 4165
rect 7935 4090 8135 4115
rect 7935 4050 7950 4090
rect 7990 4050 8070 4090
rect 8110 4050 8135 4090
rect 7935 4035 8135 4050
rect 7340 2320 10025 2350
rect 7340 2270 7415 2320
rect 7465 2270 9850 2320
rect 9900 2270 9950 2320
rect 10000 2270 10025 2320
rect 7340 2220 10025 2270
rect 7340 2170 7415 2220
rect 7465 2170 9850 2220
rect 9900 2170 9950 2220
rect 10000 2170 10025 2220
rect 7340 2150 10025 2170
rect -3145 525 645 555
rect -3145 475 -3125 525
rect -3075 475 -3025 525
rect -2975 490 645 525
rect -2975 480 465 490
rect -2975 475 -715 480
rect -3145 440 -715 475
rect -675 440 -610 480
rect -570 475 465 480
rect -570 440 -135 475
rect -3145 435 -135 440
rect -95 435 -25 475
rect 15 450 465 475
rect 505 450 585 490
rect 625 450 645 490
rect 15 435 645 450
rect -3145 425 645 435
rect -3145 375 -3125 425
rect -3075 375 -3025 425
rect -2975 410 645 425
rect -2975 375 -715 410
rect -3145 370 -715 375
rect -675 370 -610 410
rect -570 405 465 410
rect -570 370 -135 405
rect -3145 365 -135 370
rect -95 365 -25 405
rect 15 370 465 405
rect 505 370 585 410
rect 625 370 645 410
rect 15 365 645 370
rect -3145 355 645 365
rect 9255 -1195 10025 -1170
rect 9255 -1235 9325 -1195
rect 9365 -1235 9855 -1195
rect 9255 -1245 9855 -1235
rect 9905 -1245 9955 -1195
rect 10005 -1245 10025 -1195
rect 9255 -1275 10025 -1245
rect 9255 -1315 9325 -1275
rect 9365 -1295 10025 -1275
rect 9365 -1315 9855 -1295
rect 9255 -1345 9855 -1315
rect 9905 -1345 9955 -1295
rect 10005 -1345 10025 -1295
rect 9255 -1370 10025 -1345
rect -2065 -1560 1380 -1540
rect -2065 -1610 -2035 -1560
rect -1985 -1610 -1935 -1560
rect -1885 -1610 1380 -1560
rect -2065 -1660 1380 -1610
rect -2065 -1710 -2035 -1660
rect -1985 -1710 -1935 -1660
rect -1885 -1670 1380 -1660
rect -1885 -1710 1190 -1670
rect 1230 -1710 1270 -1670
rect 1310 -1710 1380 -1670
rect -2065 -1740 1380 -1710
rect 6580 -1785 10990 -1770
rect 6580 -1825 6650 -1785
rect 6690 -1790 10990 -1785
rect 6690 -1825 10815 -1790
rect 6580 -1840 10815 -1825
rect 10865 -1840 10915 -1790
rect 10965 -1840 10990 -1790
rect 6580 -1890 10990 -1840
rect 6580 -1905 10815 -1890
rect 6580 -1945 6650 -1905
rect 6690 -1940 10815 -1905
rect 10865 -1940 10915 -1890
rect 10965 -1940 10990 -1890
rect 6690 -1945 10990 -1940
rect 6580 -1970 10990 -1945
rect -3145 -2110 -960 -2095
rect -3145 -2115 -1145 -2110
rect -3145 -2165 -3120 -2115
rect -3070 -2165 -3020 -2115
rect -2970 -2150 -1145 -2115
rect -1105 -2150 -1020 -2110
rect -980 -2150 -960 -2110
rect -2970 -2165 -960 -2150
rect -3145 -2185 -960 -2165
rect -3145 -2215 -1145 -2185
rect -3145 -2265 -3120 -2215
rect -3070 -2265 -3020 -2215
rect -2970 -2225 -1145 -2215
rect -1105 -2225 -1020 -2185
rect -980 -2225 -960 -2185
rect -2970 -2265 -960 -2225
rect -3145 -2295 -960 -2265
rect -1645 -2815 1245 -2735
rect -1645 -2855 -715 -2815
rect -675 -2855 -615 -2815
rect -575 -2855 150 -2815
rect 190 -2855 250 -2815
rect 290 -2855 1070 -2815
rect 1110 -2855 1170 -2815
rect 1210 -2855 1245 -2815
rect -1645 -2885 1245 -2855
rect -1645 -2925 -715 -2885
rect -675 -2925 -615 -2885
rect -575 -2925 150 -2885
rect 190 -2925 250 -2885
rect 290 -2925 1070 -2885
rect 1110 -2925 1170 -2885
rect 1210 -2925 1245 -2885
rect -1645 -2935 1245 -2925
rect -1645 -3130 -1435 -2935
rect -1725 -3135 -1435 -3130
rect -2065 -3160 -1435 -3135
rect -2065 -3210 -2045 -3160
rect -1995 -3210 -1945 -3160
rect -1895 -3210 -1435 -3160
rect -2065 -3260 -1435 -3210
rect -2065 -3310 -2045 -3260
rect -1995 -3310 -1945 -3260
rect -1895 -3310 -1435 -3260
rect -2065 -3335 -1435 -3310
rect 9255 -3495 10025 -3470
rect -2065 -3540 -740 -3515
rect -2065 -3590 -2045 -3540
rect -1995 -3590 -1945 -3540
rect -1895 -3590 -740 -3540
rect -2065 -3605 -740 -3590
rect -2065 -3640 -965 -3605
rect -2065 -3690 -2045 -3640
rect -1995 -3690 -1945 -3640
rect -1895 -3645 -965 -3640
rect -925 -3645 -885 -3605
rect -845 -3645 -805 -3605
rect -765 -3645 -740 -3605
rect -1895 -3660 -740 -3645
rect 9255 -3535 9850 -3495
rect 9255 -3575 9325 -3535
rect 9365 -3545 9850 -3535
rect 9900 -3545 9950 -3495
rect 10000 -3545 10025 -3495
rect 9365 -3575 10025 -3545
rect 9255 -3595 10025 -3575
rect 9255 -3615 9850 -3595
rect 9255 -3655 9325 -3615
rect 9365 -3645 9850 -3615
rect 9900 -3645 9950 -3595
rect 10000 -3645 10025 -3595
rect 9365 -3655 10025 -3645
rect -1895 -3690 -1865 -3660
rect 9255 -3670 10025 -3655
rect -2065 -3715 -1865 -3690
rect 6125 -4115 6325 -4110
rect 6125 -4155 6135 -4115
rect 6175 -4155 6255 -4115
rect 6295 -4155 6325 -4115
rect 6125 -4165 6325 -4155
rect 6125 -4215 6140 -4165
rect 6190 -4215 6240 -4165
rect 6290 -4215 6325 -4165
rect 6125 -4220 6325 -4215
rect -1620 -4630 -1420 -4620
rect -1620 -4670 -1605 -4630
rect -1565 -4670 -1490 -4630
rect -1450 -4670 -1420 -4630
rect -1620 -4690 -1420 -4670
rect -1620 -4740 -1605 -4690
rect -1555 -4740 -1505 -4690
rect -1455 -4740 -1420 -4690
rect 290 -4630 490 -4620
rect 290 -4670 305 -4630
rect 345 -4670 420 -4630
rect 460 -4670 490 -4630
rect 290 -4685 490 -4670
rect 290 -4735 300 -4685
rect 350 -4735 400 -4685
rect 450 -4735 490 -4685
rect 290 -4740 490 -4735
rect -1620 -4750 -1420 -4740
rect 4000 -4845 4195 -4830
rect 4000 -4885 4020 -4845
rect 4060 -4885 4130 -4845
rect 4170 -4885 4195 -4845
rect 4000 -4900 4195 -4885
rect 4000 -4950 4015 -4900
rect 4065 -4950 4125 -4900
rect 4175 -4950 4195 -4900
rect 4000 -4955 4195 -4950
rect 8035 -4845 8230 -4830
rect 8035 -4885 8050 -4845
rect 8090 -4885 8170 -4845
rect 8210 -4885 8230 -4845
rect 8035 -4910 8230 -4885
rect 8035 -4960 8055 -4910
rect 8105 -4960 8155 -4910
rect 8205 -4960 8230 -4910
rect 8035 -4970 8230 -4960
rect -2074 -5755 10030 -5678
rect -2074 -5805 -2035 -5755
rect -1985 -5805 -1935 -5755
rect -1885 -5760 10030 -5755
rect -1885 -5805 4020 -5760
rect -2074 -5810 4020 -5805
rect 4070 -5810 4120 -5760
rect 4170 -5810 8060 -5760
rect 8110 -5810 8160 -5760
rect 8210 -5765 10030 -5760
rect 8210 -5810 9845 -5765
rect -2074 -5815 9845 -5810
rect 9895 -5815 9945 -5765
rect 9995 -5815 10030 -5765
rect -2074 -5855 10030 -5815
rect -2074 -5905 -2035 -5855
rect -1985 -5905 -1935 -5855
rect -1885 -5860 10030 -5855
rect -1885 -5905 4020 -5860
rect -2074 -5910 4020 -5905
rect 4070 -5910 4120 -5860
rect 4170 -5910 8060 -5860
rect 8110 -5910 8160 -5860
rect 8210 -5865 10030 -5860
rect 8210 -5910 9845 -5865
rect -2074 -5915 9845 -5910
rect 9895 -5915 9945 -5865
rect 9995 -5915 10030 -5865
rect -2074 -5950 10030 -5915
rect -3162 -6845 11050 -6766
rect -3162 -6860 -1600 -6845
rect -3162 -6910 -3120 -6860
rect -3070 -6910 -3020 -6860
rect -2970 -6895 -1600 -6860
rect -1550 -6895 -1500 -6845
rect -1450 -6855 11050 -6845
rect -1450 -6895 315 -6855
rect -2970 -6905 315 -6895
rect 365 -6905 415 -6855
rect 465 -6905 6150 -6855
rect 6200 -6905 6250 -6855
rect 6300 -6865 11050 -6855
rect 6300 -6905 10810 -6865
rect -2970 -6910 10810 -6905
rect -3162 -6915 10810 -6910
rect 10860 -6915 10910 -6865
rect 10960 -6915 11050 -6865
rect -3162 -6945 11050 -6915
rect -3162 -6960 -1600 -6945
rect -3162 -7010 -3120 -6960
rect -3070 -7010 -3020 -6960
rect -2970 -6995 -1600 -6960
rect -1550 -6995 -1500 -6945
rect -1450 -6955 11050 -6945
rect -1450 -6995 315 -6955
rect -2970 -7005 315 -6995
rect 365 -7005 415 -6955
rect 465 -7005 6150 -6955
rect 6200 -7005 6250 -6955
rect 6300 -6965 11050 -6955
rect 6300 -7005 10810 -6965
rect -2970 -7010 10810 -7005
rect -3162 -7015 10810 -7010
rect 10860 -7015 10910 -6965
rect 10960 -7015 11050 -6965
rect -3162 -7038 11050 -7015
rect -7645 -13150 -6935 -13085
rect -7645 -13220 -7595 -13150
rect -7525 -13220 -7455 -13150
rect -7385 -13220 -7315 -13150
rect -7245 -13220 -7175 -13150
rect -7105 -13220 -7040 -13150
rect -6970 -13220 -6935 -13150
rect -7645 -13285 -6935 -13220
<< via3 >>
rect -3120 5820 -3070 5870
rect -3020 5820 -2970 5870
rect 265 5855 315 5905
rect 365 5855 415 5905
rect 2130 5840 2180 5890
rect 2230 5840 2280 5890
rect 5540 5815 5590 5865
rect 5640 5815 5690 5865
rect 7960 5820 8010 5870
rect 8060 5820 8110 5870
rect 10810 5815 10860 5865
rect 10910 5815 10960 5865
rect -3120 5720 -3070 5770
rect -3020 5720 -2970 5770
rect 265 5755 315 5805
rect 365 5755 415 5805
rect 2130 5740 2180 5790
rect 2230 5740 2280 5790
rect 5540 5715 5590 5765
rect 5640 5715 5690 5765
rect 7960 5720 8010 5770
rect 8060 5720 8110 5770
rect 10810 5715 10860 5765
rect 10910 5715 10960 5765
rect -2035 4820 -1985 4870
rect -1935 4820 -1885 4870
rect 9850 4815 9900 4865
rect 9950 4815 10000 4865
rect -2035 4720 -1985 4770
rect -1935 4720 -1885 4770
rect 9850 4715 9900 4765
rect 9950 4715 10000 4765
rect 265 4125 315 4175
rect 365 4125 415 4175
rect 255 4090 315 4100
rect 255 4050 265 4090
rect 265 4050 305 4090
rect 305 4050 315 4090
rect 255 4040 315 4050
rect 375 4090 435 4100
rect 375 4050 385 4090
rect 385 4050 425 4090
rect 425 4050 435 4090
rect 375 4040 435 4050
rect 2130 4125 2180 4175
rect 2230 4125 2280 4175
rect 5540 4125 5590 4175
rect 5640 4125 5690 4175
rect 7950 4115 8000 4165
rect 8065 4115 8115 4165
rect 9850 2270 9900 2320
rect 9950 2270 10000 2320
rect 9850 2170 9900 2220
rect 9950 2170 10000 2220
rect -3125 475 -3075 525
rect -3025 475 -2975 525
rect -3125 375 -3075 425
rect -3025 375 -2975 425
rect 9855 -1245 9905 -1195
rect 9955 -1245 10005 -1195
rect 9855 -1345 9905 -1295
rect 9955 -1345 10005 -1295
rect -2035 -1610 -1985 -1560
rect -1935 -1610 -1885 -1560
rect -2035 -1710 -1985 -1660
rect -1935 -1710 -1885 -1660
rect 10815 -1840 10865 -1790
rect 10915 -1840 10965 -1790
rect 10815 -1940 10865 -1890
rect 10915 -1940 10965 -1890
rect -3120 -2165 -3070 -2115
rect -3020 -2165 -2970 -2115
rect -3120 -2265 -3070 -2215
rect -3020 -2265 -2970 -2215
rect -2045 -3210 -1995 -3160
rect -1945 -3210 -1895 -3160
rect -2045 -3310 -1995 -3260
rect -1945 -3310 -1895 -3260
rect -2045 -3590 -1995 -3540
rect -1945 -3590 -1895 -3540
rect -2045 -3690 -1995 -3640
rect -1945 -3690 -1895 -3640
rect 9850 -3545 9900 -3495
rect 9950 -3545 10000 -3495
rect 9850 -3645 9900 -3595
rect 9950 -3645 10000 -3595
rect 6140 -4215 6190 -4165
rect 6240 -4215 6290 -4165
rect -1605 -4740 -1555 -4690
rect -1505 -4740 -1455 -4690
rect 300 -4735 350 -4685
rect 400 -4735 450 -4685
rect 4015 -4950 4065 -4900
rect 4125 -4950 4175 -4900
rect 8055 -4960 8105 -4910
rect 8155 -4960 8205 -4910
rect -2035 -5805 -1985 -5755
rect -1935 -5805 -1885 -5755
rect 4020 -5810 4070 -5760
rect 4120 -5810 4170 -5760
rect 8060 -5810 8110 -5760
rect 8160 -5810 8210 -5760
rect 9845 -5815 9895 -5765
rect 9945 -5815 9995 -5765
rect -2035 -5905 -1985 -5855
rect -1935 -5905 -1885 -5855
rect 4020 -5910 4070 -5860
rect 4120 -5910 4170 -5860
rect 8060 -5910 8110 -5860
rect 8160 -5910 8210 -5860
rect 9845 -5915 9895 -5865
rect 9945 -5915 9995 -5865
rect -3120 -6910 -3070 -6860
rect -3020 -6910 -2970 -6860
rect -1600 -6895 -1550 -6845
rect -1500 -6895 -1450 -6845
rect 315 -6905 365 -6855
rect 415 -6905 465 -6855
rect 6150 -6905 6200 -6855
rect 6250 -6905 6300 -6855
rect 10810 -6915 10860 -6865
rect 10910 -6915 10960 -6865
rect -3120 -7010 -3070 -6960
rect -3020 -7010 -2970 -6960
rect -1600 -6995 -1550 -6945
rect -1500 -6995 -1450 -6945
rect 315 -7005 365 -6955
rect 415 -7005 465 -6955
rect 6150 -7005 6200 -6955
rect 6250 -7005 6300 -6955
rect 10810 -7015 10860 -6965
rect 10910 -7015 10960 -6965
<< metal4 >>
rect -3162 5870 -2890 5950
rect -3162 5820 -3120 5870
rect -3070 5820 -3020 5870
rect -2970 5820 -2890 5870
rect -3162 5770 -2890 5820
rect -3162 5720 -3120 5770
rect -3070 5720 -3020 5770
rect -2970 5720 -2890 5770
rect -3162 525 -2890 5720
rect 245 5905 445 5950
rect 245 5855 265 5905
rect 315 5855 365 5905
rect 415 5855 445 5905
rect 245 5805 445 5855
rect 245 5755 265 5805
rect 315 5755 365 5805
rect 415 5755 445 5805
rect -3162 475 -3125 525
rect -3075 475 -3025 525
rect -2975 475 -2890 525
rect -3162 425 -2890 475
rect -3162 375 -3125 425
rect -3075 375 -3025 425
rect -2975 375 -2890 425
rect -3162 -2115 -2890 375
rect -3162 -2165 -3120 -2115
rect -3070 -2165 -3020 -2115
rect -2970 -2165 -2890 -2115
rect -3162 -2215 -2890 -2165
rect -3162 -2265 -3120 -2215
rect -3070 -2265 -3020 -2215
rect -2970 -2265 -2890 -2215
rect -3162 -6860 -2890 -2265
rect -2074 4870 -1802 4930
rect -2074 4820 -2035 4870
rect -1985 4820 -1935 4870
rect -1885 4820 -1802 4870
rect -2074 4770 -1802 4820
rect -2074 4720 -2035 4770
rect -1985 4720 -1935 4770
rect -1885 4720 -1802 4770
rect -2074 -1560 -1802 4720
rect 245 4175 445 5755
rect 245 4125 265 4175
rect 315 4125 365 4175
rect 415 4125 445 4175
rect 245 4100 445 4125
rect 245 4040 255 4100
rect 315 4040 375 4100
rect 435 4040 445 4100
rect 245 3995 445 4040
rect 2110 5890 2310 5950
rect 2110 5840 2130 5890
rect 2180 5840 2230 5890
rect 2280 5840 2310 5890
rect 2110 5790 2310 5840
rect 2110 5740 2130 5790
rect 2180 5740 2230 5790
rect 2280 5740 2310 5790
rect 2110 4175 2310 5740
rect 2110 4125 2130 4175
rect 2180 4125 2230 4175
rect 2280 4125 2310 4175
rect 2110 3995 2310 4125
rect 5520 5865 5720 5895
rect 5520 5815 5540 5865
rect 5590 5815 5640 5865
rect 5690 5815 5720 5865
rect 5520 5765 5720 5815
rect 5520 5715 5540 5765
rect 5590 5715 5640 5765
rect 5690 5715 5720 5765
rect 5520 4175 5720 5715
rect 5520 4125 5540 4175
rect 5590 4125 5640 4175
rect 5690 4125 5720 4175
rect 5520 3995 5720 4125
rect 7935 5870 8135 5895
rect 7935 5820 7960 5870
rect 8010 5820 8060 5870
rect 8110 5820 8135 5870
rect 7935 5770 8135 5820
rect 7935 5720 7960 5770
rect 8010 5720 8060 5770
rect 8110 5720 8135 5770
rect 7935 4165 8135 5720
rect 10778 5865 11050 5950
rect 10778 5815 10810 5865
rect 10860 5815 10910 5865
rect 10960 5815 11050 5865
rect 10778 5765 11050 5815
rect 10778 5715 10810 5765
rect 10860 5715 10910 5765
rect 10960 5715 11050 5765
rect 7935 4115 7950 4165
rect 8000 4115 8065 4165
rect 8115 4115 8135 4165
rect 7935 3995 8135 4115
rect 9758 4865 10030 4930
rect 9758 4815 9850 4865
rect 9900 4815 9950 4865
rect 10000 4815 10030 4865
rect 9758 4765 10030 4815
rect 9758 4715 9850 4765
rect 9900 4715 9950 4765
rect 10000 4715 10030 4765
rect -2074 -1610 -2035 -1560
rect -1985 -1610 -1935 -1560
rect -1885 -1610 -1802 -1560
rect -2074 -1660 -1802 -1610
rect -2074 -1710 -2035 -1660
rect -1985 -1710 -1935 -1660
rect -1885 -1710 -1802 -1660
rect -2074 -3160 -1802 -1710
rect -2074 -3210 -2045 -3160
rect -1995 -3210 -1945 -3160
rect -1895 -3210 -1802 -3160
rect -2074 -3260 -1802 -3210
rect -2074 -3310 -2045 -3260
rect -1995 -3310 -1945 -3260
rect -1895 -3310 -1802 -3260
rect -2074 -3540 -1802 -3310
rect -2074 -3590 -2045 -3540
rect -1995 -3590 -1945 -3540
rect -1895 -3590 -1802 -3540
rect -2074 -3640 -1802 -3590
rect -2074 -3690 -2045 -3640
rect -1995 -3690 -1945 -3640
rect -1895 -3690 -1802 -3640
rect -2074 -5755 -1802 -3690
rect 9758 2320 10030 4715
rect 9758 2270 9850 2320
rect 9900 2270 9950 2320
rect 10000 2270 10030 2320
rect 9758 2220 10030 2270
rect 9758 2170 9850 2220
rect 9900 2170 9950 2220
rect 10000 2170 10030 2220
rect 9758 -1195 10030 2170
rect 9758 -1245 9855 -1195
rect 9905 -1245 9955 -1195
rect 10005 -1245 10030 -1195
rect 9758 -1295 10030 -1245
rect 9758 -1345 9855 -1295
rect 9905 -1345 9955 -1295
rect 10005 -1345 10030 -1295
rect 9758 -3495 10030 -1345
rect 9758 -3545 9850 -3495
rect 9900 -3545 9950 -3495
rect 10000 -3545 10030 -3495
rect 9758 -3595 10030 -3545
rect 9758 -3645 9850 -3595
rect 9900 -3645 9950 -3595
rect 10000 -3645 10030 -3595
rect 6125 -4165 6325 -4060
rect 6125 -4215 6140 -4165
rect 6190 -4215 6240 -4165
rect 6290 -4215 6325 -4165
rect -2074 -5805 -2035 -5755
rect -1985 -5805 -1935 -5755
rect -1885 -5805 -1802 -5755
rect -2074 -5855 -1802 -5805
rect -2074 -5905 -2035 -5855
rect -1985 -5905 -1935 -5855
rect -1885 -5905 -1802 -5855
rect -2074 -5950 -1802 -5905
rect -1620 -4690 -1420 -4575
rect -1620 -4740 -1605 -4690
rect -1555 -4740 -1505 -4690
rect -1455 -4740 -1420 -4690
rect -3162 -6910 -3120 -6860
rect -3070 -6910 -3020 -6860
rect -2970 -6910 -2890 -6860
rect -3162 -6960 -2890 -6910
rect -3162 -7010 -3120 -6960
rect -3070 -7010 -3020 -6960
rect -2970 -7010 -2890 -6960
rect -3162 -7038 -2890 -7010
rect -1620 -6845 -1420 -4740
rect -1620 -6895 -1600 -6845
rect -1550 -6895 -1500 -6845
rect -1450 -6895 -1420 -6845
rect -1620 -6945 -1420 -6895
rect -1620 -6995 -1600 -6945
rect -1550 -6995 -1500 -6945
rect -1450 -6995 -1420 -6945
rect -1620 -7040 -1420 -6995
rect 290 -4685 490 -4570
rect 290 -4735 300 -4685
rect 350 -4735 400 -4685
rect 450 -4735 490 -4685
rect 290 -6855 490 -4735
rect 4000 -4900 4195 -4775
rect 4000 -4950 4015 -4900
rect 4065 -4950 4125 -4900
rect 4175 -4950 4195 -4900
rect 4000 -5760 4195 -4950
rect 4000 -5810 4020 -5760
rect 4070 -5810 4120 -5760
rect 4170 -5810 4195 -5760
rect 4000 -5860 4195 -5810
rect 4000 -5910 4020 -5860
rect 4070 -5910 4120 -5860
rect 4170 -5910 4195 -5860
rect 4000 -5935 4195 -5910
rect 290 -6905 315 -6855
rect 365 -6905 415 -6855
rect 465 -6905 490 -6855
rect 290 -6955 490 -6905
rect 290 -7005 315 -6955
rect 365 -7005 415 -6955
rect 465 -7005 490 -6955
rect 290 -7035 490 -7005
rect 6125 -6855 6325 -4215
rect 8035 -4910 8230 -4780
rect 8035 -4960 8055 -4910
rect 8105 -4960 8155 -4910
rect 8205 -4960 8230 -4910
rect 8035 -5760 8230 -4960
rect 8035 -5810 8060 -5760
rect 8110 -5810 8160 -5760
rect 8210 -5810 8230 -5760
rect 8035 -5860 8230 -5810
rect 8035 -5910 8060 -5860
rect 8110 -5910 8160 -5860
rect 8210 -5910 8230 -5860
rect 8035 -5935 8230 -5910
rect 9758 -5765 10030 -3645
rect 9758 -5815 9845 -5765
rect 9895 -5815 9945 -5765
rect 9995 -5815 10030 -5765
rect 9758 -5865 10030 -5815
rect 9758 -5915 9845 -5865
rect 9895 -5915 9945 -5865
rect 9995 -5915 10030 -5865
rect 9758 -5950 10030 -5915
rect 10778 -1790 11050 5715
rect 10778 -1840 10815 -1790
rect 10865 -1840 10915 -1790
rect 10965 -1840 11050 -1790
rect 10778 -1890 11050 -1840
rect 10778 -1940 10815 -1890
rect 10865 -1940 10915 -1890
rect 10965 -1940 11050 -1890
rect 6125 -6905 6150 -6855
rect 6200 -6905 6250 -6855
rect 6300 -6905 6325 -6855
rect 6125 -6955 6325 -6905
rect 6125 -7005 6150 -6955
rect 6200 -7005 6250 -6955
rect 6300 -7005 6325 -6955
rect 6125 -7035 6325 -7005
rect 10778 -6865 11050 -1940
rect 10778 -6915 10810 -6865
rect 10860 -6915 10910 -6865
rect 10960 -6915 11050 -6865
rect 10778 -6965 11050 -6915
rect 10778 -7015 10810 -6965
rect 10860 -7015 10910 -6965
rect 10960 -7015 11050 -6965
rect 10778 -7038 11050 -7015
use ALib_DCO  ALib_DCO_0 ./../dco
timestamp 1730531556
transform 1 0 2600 0 1 -2595
box 500 -2235 6705 2990
use ALib_VCO  ALib_VCO_0 ./../vco
timestamp 1730639796
transform 1 0 -1010 0 1 520
box 0 140 10320 3515
use DLib_Quantizer  DLib_Quantizer_0 ./../quantizer
timestamp 1730532965
transform 1 0 -1105 0 1 -2315
box 95 -355 2945 365
use DLib_UpDownCounter  DLib_UpDownCounter_0 ./../count
timestamp 1730536752
transform 1 0 -570 0 1 -2993
box -440 -1577 1570 -220
use DLib_UpDownCounter  DLib_UpDownCounter_1
timestamp 1730536752
transform 1 0 -570 0 1 172
box -440 -1577 1570 -220
<< labels >>
flabel metal3 -2970 5678 -535 5950 1 FreeSans 1088 0 0 0 VDDA
port 7 nsew power input
flabel metal3 8194 4658 9758 4930 1 FreeSans 1088 0 0 0 GND
port 8 nsew ground input
rlabel locali 365 4035 365 4035 1 VDDA
port 4 n
<< end >>
