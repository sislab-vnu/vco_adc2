* NGSPICE file created from mag_vco_aux_inv.ext - technology: sky130A

.subckt mag_vco_aux_inv A VPWR VGND Y VCCA GND
X0 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

