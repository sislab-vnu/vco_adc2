* NGSPICE file created from obr.ext - technology: sky130A

.subckt p_br1 G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
.ends

.subckt p_br2 G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
.ends

.subckt obr s_1 g_1 d_1 s_2 g_2 d_2
Xp_br1_0 g_1 s_1 d_1 s_1 p_br1
Xp_br2_0 g_2 s_2 d_2 s_2 p_br2
.ends

