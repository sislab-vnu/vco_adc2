VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc2
  CLASS BLOCK ;
  FOREIGN vco_adc2 ;
  ORIGIN 77.180 133.620 ;
  SIZE 285.330 BY 295.770 ;
  PIN vbias_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met3 ;
        RECT -77.180 127.500 -69.020 132.260 ;
    END
  END vbias_12
  PIN vbias_34
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER met3 ;
        RECT -77.180 -133.620 -69.020 -128.860 ;
    END
  END vbias_34
  PIN analog_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.570 160.310 208.150 162.150 ;
    END
  END analog_in
  PIN enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.437000 ;
    PORT
      LAYER met2 ;
        RECT -6.240 -133.170 -3.480 -126.270 ;
    END
  END enable_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER met2 ;
        RECT -37.030 -133.170 -34.730 -126.270 ;
    END
  END clk
  PIN quantizer_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 14.000 -133.150 16.760 -125.790 ;
    END
  END quantizer_out
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -44.540 -117.300 -41.820 59.500 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.540 -117.300 124.780 -114.580 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.540 56.780 124.780 59.500 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -20.740 -95.540 -18.020 49.300 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.740 -95.540 100.300 -92.820 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.740 46.580 100.300 49.300 ;
    END
  END vssa1
  OBS
      LAYER li1 ;
        RECT -14.000 -50.500 93.100 40.350 ;
      LAYER met1 ;
        RECT -14.000 -50.500 93.050 40.350 ;
      LAYER met2 ;
        RECT -77.180 160.030 197.290 160.310 ;
        RECT -77.180 -125.510 199.450 160.030 ;
        RECT -77.180 -125.990 13.720 -125.510 ;
        RECT -77.180 -133.450 -37.310 -125.990 ;
        RECT -34.450 -133.450 -6.520 -125.990 ;
        RECT -3.200 -133.430 13.720 -125.990 ;
        RECT 17.040 -133.430 199.450 -125.510 ;
        RECT -3.200 -133.450 199.450 -133.430 ;
        RECT -77.180 -133.620 199.450 -133.450 ;
      LAYER met3 ;
        RECT -44.650 49.700 124.800 56.380 ;
        RECT -44.650 46.180 -21.140 49.700 ;
        RECT 100.700 46.180 124.800 49.700 ;
        RECT -44.650 -92.420 124.800 46.180 ;
        RECT -44.650 -95.940 -21.140 -92.420 ;
        RECT 100.700 -95.940 124.800 -92.420 ;
        RECT -44.650 -114.180 124.800 -95.940 ;
      LAYER met4 ;
        RECT -41.420 49.700 124.800 59.800 ;
        RECT -41.420 -95.940 -21.140 49.700 ;
        RECT -17.620 -95.940 124.800 49.700 ;
        RECT -41.420 -117.400 124.800 -95.940 ;
  END
END vco_adc2
END LIBRARY

