* NGSPICE file created from DLib_Quantizer.ext - technology: sky130A






.subckt DLib_Quantizer D CLK Dout FBack VDDA GND
Xsky130_fd_sc_hd__dlygate4sd3_1_0 CLK GND GND VDDA VDDA DL1 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_1 DL1 GND GND VDDA VDDA DL2 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__inv_2_0 FBack_inv GND GND VDDA VDDA FBack sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_0 D GND GND VDDA VDDA sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dlygate4sd3_1_2 DL2 GND GND VDDA VDDA DL3 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_3 DL3 GND GND VDDA VDDA DL4 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_4 DL4 GND GND VDDA VDDA DL5 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_5 DL5 GND GND VDDA VDDA CLK_dly sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__nand2_1_0 CLK_dly Dout GND GND VDDA VDDA FBack_inv sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_0 CLK sky130_fd_sc_hd__buf_2_0/X GND GND VDDA VDDA Dout
+ sky130_fd_sc_hd__dfxtp_1
.ends


