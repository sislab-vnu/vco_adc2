* NGSPICE file created from save.ext - technology: sky130A

.subckt save A VPWR VGND Y
X0 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
X1 Y A VPWR w_n130_n80# sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
.ends

