* NGSPICE file created from vco_main_inv.ext - technology: sky130A

.subckt vco_main_inv A VPWR VGND Y VCCA GND
X0 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends


