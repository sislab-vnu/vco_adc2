magic
tech sky130A
timestamp 1725875793
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 0 0 1 0
box -19 -24 249 296
<< properties >>
string FIXED_BBOX 1
<< end >>
