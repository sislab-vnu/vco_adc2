magic
tech sky130A
magscale 1 2
timestamp 1723880701
<< nwell >>
rect -344 -766 -28 -450
rect 1942 -750 2258 -450
rect -298 -770 -46 -766
rect 1942 -772 2404 -750
rect 1968 -774 2404 -772
rect -868 -1814 -698 -1492
rect 1586 -1908 1814 -1586
rect -192 -2824 -22 -2822
rect 1914 -2824 2130 -2822
rect -192 -3144 -42 -2824
rect 1914 -2828 2056 -2824
rect 1958 -3144 2056 -2828
<< pwell >>
rect 1830 -876 2398 -830
rect -332 -1010 -4 -876
rect 1830 -982 2310 -876
rect 2314 -878 2398 -876
rect 2320 -880 2398 -878
rect 2326 -982 2398 -880
rect 1830 -1012 2398 -982
rect -868 -2056 -664 -1872
rect 1568 -2010 1854 -1964
rect 1568 -2148 1860 -2010
rect -228 -2766 70 -2582
rect 1924 -2720 2096 -2582
<< psubdiff >>
rect 2172 -902 2230 -870
rect 2172 -936 2184 -902
rect 2218 -936 2230 -902
rect 2172 -970 2230 -936
rect -810 -1942 -752 -1908
rect -810 -1976 -798 -1942
rect -764 -1976 -752 -1942
rect -810 -2008 -752 -1976
rect 1678 -2050 1736 -2014
rect 1678 -2084 1690 -2050
rect 1724 -2084 1736 -2050
rect 1678 -2114 1736 -2084
rect 1974 -2636 2032 -2602
rect 1974 -2670 1986 -2636
rect 2020 -2670 2032 -2636
rect 1974 -2702 2032 -2670
<< nsubdiff >>
rect 2058 -602 2116 -568
rect 2058 -638 2070 -602
rect 2104 -638 2116 -602
rect 2058 -668 2116 -638
rect -810 -1656 -752 -1626
rect -810 -1690 -798 -1656
rect -764 -1690 -752 -1656
rect -810 -1726 -752 -1690
rect 1676 -1704 1734 -1668
rect 1676 -1738 1688 -1704
rect 1722 -1738 1734 -1704
rect 1676 -1768 1734 -1738
rect 1976 -2958 2034 -2924
rect 1976 -2992 1986 -2958
rect 2020 -2992 2034 -2958
rect 1976 -3022 2034 -2992
<< psubdiffcont >>
rect 2184 -936 2218 -902
rect -798 -1976 -764 -1942
rect 1690 -2084 1724 -2050
rect 1986 -2670 2020 -2636
<< nsubdiffcont >>
rect 2070 -638 2104 -602
rect -798 -1690 -764 -1656
rect 1688 -1738 1722 -1704
rect 1986 -2992 2020 -2958
<< locali >>
rect 2058 -602 2116 -568
rect 2058 -638 2070 -602
rect 2104 -638 2116 -602
rect 2058 -668 2116 -638
rect 2172 -902 2230 -870
rect 2172 -936 2184 -902
rect 2218 -936 2230 -902
rect 2172 -970 2230 -936
rect -810 -1656 -752 -1626
rect -810 -1690 -798 -1656
rect -764 -1690 -752 -1656
rect -810 -1726 -752 -1690
rect 1676 -1704 1734 -1668
rect 1676 -1738 1688 -1704
rect 1722 -1738 1734 -1704
rect 1676 -1768 1734 -1738
rect 1532 -1894 1736 -1818
rect 1664 -1898 1736 -1894
rect -810 -1942 -752 -1908
rect -810 -1976 -798 -1942
rect -764 -1976 -752 -1942
rect 1664 -1972 1866 -1898
rect -810 -2008 -752 -1976
rect 1678 -2050 1736 -2014
rect 1678 -2084 1690 -2050
rect 1724 -2084 1736 -2050
rect 1678 -2114 1736 -2084
rect 1974 -2636 2032 -2602
rect 1974 -2670 1986 -2636
rect 2020 -2670 2032 -2636
rect 1974 -2702 2032 -2670
rect 1976 -2958 2034 -2924
rect 1976 -2992 1986 -2958
rect 2020 -2992 2034 -2958
rect 1976 -3022 2034 -2992
<< viali >>
rect 2070 -638 2104 -602
rect -482 -684 -448 -650
rect 2494 -686 2528 -652
rect -660 -816 -626 -782
rect 18 -802 52 -768
rect 340 -800 374 -766
rect 1792 -818 1826 -784
rect 2316 -818 2350 -784
rect 2184 -936 2218 -902
rect -798 -1690 -764 -1656
rect -552 -1692 -518 -1658
rect 1688 -1738 1722 -1704
rect -634 -1858 -600 -1824
rect -798 -1976 -764 -1942
rect 1016 -1952 1050 -1918
rect 1132 -1954 1166 -1920
rect 1690 -2084 1724 -2050
rect 1986 -2670 2020 -2636
rect -296 -2812 -262 -2778
rect 86 -2810 120 -2776
rect 1538 -2818 1572 -2784
rect 1860 -2826 1894 -2792
rect 2388 -2810 2422 -2776
rect -380 -2980 -346 -2946
rect 2212 -2942 2246 -2908
rect 1986 -2992 2020 -2958
<< metal1 >>
rect -492 -608 -432 -562
rect 2058 -602 2116 -568
rect -492 -650 -96 -608
rect -492 -684 -482 -650
rect -448 -668 -96 -650
rect 2058 -638 2070 -602
rect 2104 -638 2116 -602
rect 2058 -668 2116 -638
rect 2486 -600 2544 -594
rect 2486 -618 2934 -600
rect 2486 -652 2864 -618
rect -448 -684 -432 -668
rect -492 -706 -432 -684
rect -736 -782 -608 -758
rect -736 -816 -660 -782
rect -626 -816 -608 -782
rect -736 -832 -608 -816
rect -156 -772 -96 -668
rect 2486 -686 2494 -652
rect 2528 -670 2864 -652
rect 2916 -670 2934 -618
rect 2528 -686 2934 -670
rect 2486 -694 2934 -686
rect 4 -768 74 -706
rect 4 -772 18 -768
rect -156 -802 18 -772
rect 52 -802 74 -768
rect -156 -832 74 -802
rect 322 -756 406 -708
rect 2486 -720 2544 -694
rect 322 -808 340 -756
rect 392 -808 406 -756
rect 2296 -772 2368 -760
rect 322 -814 406 -808
rect 1786 -784 2368 -772
rect 4 -836 74 -832
rect 1786 -818 1792 -784
rect 1826 -818 2316 -784
rect 2350 -818 2368 -784
rect 1786 -834 2368 -818
rect 702 -842 804 -836
rect 702 -894 720 -842
rect 772 -894 804 -842
rect 702 -924 804 -894
rect 2010 -1074 2090 -834
rect 2303 -836 2368 -834
rect 2172 -902 2230 -870
rect 2172 -936 2184 -902
rect 2218 -936 2230 -902
rect 2172 -970 2230 -936
rect -312 -1288 804 -1282
rect -312 -1340 724 -1288
rect 776 -1340 804 -1288
rect -312 -1346 804 -1340
rect -810 -1656 -752 -1626
rect -810 -1690 -798 -1656
rect -764 -1690 -752 -1656
rect -810 -1726 -752 -1690
rect -568 -1640 -498 -1630
rect -312 -1640 -252 -1346
rect 2008 -1420 2092 -1074
rect -568 -1658 -252 -1640
rect -568 -1692 -552 -1658
rect -518 -1692 -252 -1658
rect -568 -1700 -252 -1692
rect 496 -1484 2092 -1420
rect -568 -1720 -498 -1700
rect -831 -1824 -584 -1808
rect -831 -1858 -634 -1824
rect -600 -1858 -584 -1824
rect -831 -1874 -584 -1858
rect 496 -1904 560 -1484
rect 1676 -1704 1734 -1668
rect 1676 -1738 1688 -1704
rect 1722 -1738 1734 -1704
rect 1676 -1768 1734 -1738
rect -810 -1942 -752 -1908
rect -810 -1976 -798 -1942
rect -764 -1976 -752 -1942
rect 496 -1918 1064 -1904
rect 496 -1952 1016 -1918
rect 1050 -1952 1064 -1918
rect 496 -1968 1064 -1952
rect 1126 -1920 1190 -1908
rect 1126 -1954 1132 -1920
rect 1166 -1954 1190 -1920
rect -810 -2008 -752 -1976
rect 1126 -2012 1190 -1954
rect -152 -2072 1190 -2012
rect 1678 -2050 1736 -2014
rect -152 -2760 -84 -2072
rect 1678 -2084 1690 -2050
rect 1724 -2084 1736 -2050
rect 1678 -2114 1736 -2084
rect 1974 -2636 2032 -2602
rect 1110 -2692 1206 -2662
rect 1110 -2744 1132 -2692
rect 1184 -2744 1206 -2692
rect 1974 -2670 1986 -2636
rect 2020 -2670 2032 -2636
rect 1974 -2702 2032 -2670
rect 1110 -2756 1206 -2744
rect -310 -2776 126 -2760
rect -310 -2778 86 -2776
rect -310 -2812 -296 -2778
rect -262 -2810 86 -2778
rect 120 -2810 126 -2776
rect -262 -2812 126 -2810
rect -310 -2828 126 -2812
rect 1490 -2784 1594 -2778
rect 1490 -2798 1538 -2784
rect 1490 -2850 1510 -2798
rect 1572 -2818 1594 -2784
rect 1562 -2850 1594 -2818
rect 1490 -2886 1594 -2850
rect 1838 -2792 1908 -2756
rect 1838 -2826 1860 -2792
rect 1894 -2794 1908 -2792
rect 2372 -2776 2558 -2758
rect 1894 -2826 2250 -2794
rect 1838 -2854 2250 -2826
rect 2372 -2810 2388 -2776
rect 2422 -2810 2558 -2776
rect 2372 -2834 2558 -2810
rect 1838 -2888 1908 -2854
rect 2198 -2874 2250 -2854
rect 2198 -2908 2252 -2874
rect -396 -2932 -328 -2908
rect -640 -2936 -328 -2932
rect -640 -2988 -626 -2936
rect -574 -2946 -328 -2936
rect -574 -2980 -380 -2946
rect -346 -2980 -328 -2946
rect -574 -2988 -328 -2980
rect -640 -2992 -328 -2988
rect -396 -3000 -328 -2992
rect 1976 -2958 2034 -2924
rect 1976 -2992 1986 -2958
rect 2020 -2992 2034 -2958
rect 2198 -2942 2212 -2908
rect 2246 -2942 2252 -2908
rect 2198 -2970 2252 -2942
rect 1976 -3022 2034 -2992
<< via1 >>
rect 2864 -670 2916 -618
rect 340 -766 392 -756
rect 340 -800 374 -766
rect 374 -800 392 -766
rect 340 -808 392 -800
rect 720 -894 772 -842
rect 724 -1340 776 -1288
rect 1132 -2744 1184 -2692
rect 1510 -2818 1538 -2798
rect 1538 -2818 1562 -2798
rect 1510 -2850 1562 -2818
rect -626 -2988 -574 -2936
<< metal2 >>
rect 2843 -618 2933 -600
rect 2843 -670 2864 -618
rect 2916 -670 2933 -618
rect 330 -756 422 -708
rect 330 -808 340 -756
rect 392 -808 422 -756
rect 330 -2314 422 -808
rect -640 -2406 422 -2314
rect 702 -842 804 -814
rect 702 -894 720 -842
rect 772 -894 804 -842
rect 702 -1288 804 -894
rect 702 -1340 724 -1288
rect 776 -1340 804 -1288
rect 702 -2320 804 -1340
rect 2843 -2278 2933 -670
rect 702 -2406 1206 -2320
rect -640 -2936 -548 -2406
rect 1110 -2692 1206 -2406
rect 1110 -2744 1132 -2692
rect 1184 -2744 1206 -2692
rect 1110 -2760 1206 -2744
rect 1490 -2368 2933 -2278
rect 1490 -2798 1580 -2368
rect 1490 -2850 1510 -2798
rect 1562 -2850 1580 -2798
rect 1490 -2886 1580 -2850
rect -640 -2988 -626 -2936
rect -574 -2988 -548 -2936
rect -640 -2992 -548 -2988
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -696 0 1 -1030
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1701704242
transform -1 0 2460 0 -1 -2562
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1701704242
transform 1 0 1846 0 1 -2168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1701704242
transform 1 0 2280 0 1 -1032
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -14 0 1 -1032
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_1
timestamp 1701704242
transform -1 0 1926 0 -1 -2562
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -672 0 1 -2074
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1701704242
transform -1 0 -224 0 -1 -2562
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 930 0 1 -2168
box -38 -48 682 592
<< end >>
