** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/ALib_IDAC.sch
.subckt ALib_IDAC Vbs1 Vbs2 Vbs3 Vbs4 Dctrl Isup VDDA GND
*.PININFO Vbs3:I Vbs4:I Vbs1:I Vbs2:I Isup:O Dctrl:I GND:I VDDA:I
x1 open GND GND VDDA VDDA lock sky130_fd_sc_hd__inv_2
XM1 net1 Vbs1 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt L=0.5 W=1.8 nf=1 m=1
XM2 Isup Vbs2 net1 net1 sky130_fd_pr__pfet_01v8_hvt L=0.5 W=1.8 nf=1 m=1
x2 Dctrl GND GND VDDA VDDA open sky130_fd_sc_hd__buf_2
XM3 net2 Vbs3 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt L=0.5 W=5.4 nf=3 m=1
XM4 add_pwr Vbs4 net2 net2 sky130_fd_pr__pfet_01v8_hvt L=0.5 W=5.4 nf=3 m=1
XM5 Isup lock add_pwr add_pwr sky130_fd_pr__pfet_01v8_hvt L=0.5 W=8 nf=2 m=1
XM6 add_pwr open Isup GND sky130_fd_pr__nfet_01v8 L=0.5 W=4 nf=2 m=1
XM7 input_R open add_pwr add_pwr sky130_fd_pr__pfet_01v8_hvt L=0.5 W=8 nf=2 m=1
XM8 add_pwr lock input_R GND sky130_fd_pr__nfet_01v8 L=0.5 W=4 nf=2 m=1
XR2 GND input_R GND sky130_fd_pr__res_xhigh_po_0p35 L=8.562 mult=1 m=1
.ends
.end
