* NGSPICE file created from DLib_freqDiv2.ext - technology: sky130A





.subckt DLib_freqDiv2 clk clkDiv2 VDDA GND
Xsky130_fd_sc_hd__buf_4_0 Q_N GND GND VDDA VDDA Q_N_buf sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_4_0 clk GND GND VDDA VDDA clkinv sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__dfxtp_1_0 clkinv Q_N_buf GND GND VDDA VDDA D sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxbp_2_0 clk D GND GND VDDA VDDA clkDiv2 Q_N sky130_fd_sc_hd__dfxbp_2
.ends


