magic
tech sky130A
timestamp 1726656757
<< poly >>
rect 500 260 730 300
rect 130 220 180 260
<< locali >>
rect 20 470 130 520
rect 20 225 60 470
rect 90 220 130 470
rect 390 470 500 520
rect 390 225 430 470
rect 180 40 220 220
rect 460 210 500 470
<< metal1 >>
rect 730 40 770 120
use p_br1  p_br1_0
timestamp 1726647752
transform 1 0 130 0 1 40
box -130 -40 108 220
use p_br2  p_br2_0
timestamp 1726647805
transform 1 0 500 0 1 40
box -130 -40 290 260
<< labels >>
rlabel locali 80 520 80 520 1 s_1
port 1 n
rlabel poly 155 260 155 260 1 g_1
port 2 n
rlabel locali 205 220 205 220 1 d_1
port 3 n
rlabel locali 445 520 445 520 1 s_2
port 4 n
rlabel poly 615 300 615 300 1 g_2
port 5 n
rlabel metal1 750 40 750 40 5 d_2
port 6 s
<< end >>
