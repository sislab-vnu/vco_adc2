magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect 1920 1260 1960 1300
rect 1920 1180 1960 1220
<< pwell >>
rect 2474 414 2566 586
<< ndiff >>
rect 2500 557 2540 560
rect 2500 523 2503 557
rect 2537 523 2540 557
rect 2500 520 2540 523
rect 2500 477 2540 480
rect 2500 443 2503 477
rect 2537 443 2540 477
rect 2500 440 2540 443
<< pdiff >>
rect 1920 1297 1960 1300
rect 1920 1263 1923 1297
rect 1957 1263 1960 1297
rect 1920 1260 1960 1263
rect 1920 1217 1960 1220
rect 1920 1183 1923 1217
rect 1957 1183 1960 1217
rect 1920 1180 1960 1183
<< ndiffc >>
rect 2503 523 2537 557
rect 2503 443 2537 477
<< pdiffc >>
rect 1923 1263 1957 1297
rect 1923 1183 1957 1217
<< poly >>
rect 1190 787 1230 790
rect 1190 753 1193 787
rect 1227 753 1230 787
rect 1190 750 1230 753
rect 1770 787 1810 790
rect 1770 753 1773 787
rect 1807 753 1810 787
rect 1770 750 1810 753
<< polycont >>
rect 1193 753 1227 787
rect 1773 753 1807 787
<< locali >>
rect 670 1660 2310 1740
rect 1040 1480 1120 1660
rect 1620 1480 1700 1660
rect 480 1297 520 1300
rect 480 1263 483 1297
rect 517 1263 520 1297
rect 480 1260 520 1263
rect 1920 1297 1960 1300
rect 1920 1263 1923 1297
rect 1957 1263 1960 1297
rect 1920 1260 1960 1263
rect 480 1217 520 1220
rect 480 1183 483 1217
rect 517 1183 520 1217
rect 480 1180 520 1183
rect 1920 1217 1960 1220
rect 1920 1183 1923 1217
rect 1957 1183 1960 1217
rect 1920 1180 1960 1183
rect 1920 1137 1960 1140
rect 1920 1103 1923 1137
rect 1957 1103 1960 1137
rect 1920 1100 1960 1103
rect 1340 977 1380 980
rect 1340 943 1343 977
rect 1377 943 1380 977
rect 1340 940 1380 943
rect 2500 977 2540 980
rect 2500 943 2503 977
rect 2537 943 2540 977
rect 2500 940 2540 943
rect 1170 787 1250 810
rect 1170 753 1193 787
rect 1227 753 1250 787
rect 1170 730 1250 753
rect 1400 787 1830 810
rect 1400 753 1773 787
rect 1807 753 1830 787
rect 1400 730 1830 753
rect 2500 557 2540 560
rect 2500 523 2503 557
rect 2537 523 2540 557
rect 2500 520 2540 523
rect 2500 477 2540 480
rect 2500 443 2503 477
rect 2537 443 2540 477
rect 2500 440 2540 443
rect 2500 397 2540 400
rect 2500 363 2503 397
rect 2537 363 2540 397
rect 2500 360 2540 363
rect 1040 80 1120 260
rect 1620 80 1700 260
rect 600 0 2220 80
<< viali >>
rect 483 1263 517 1297
rect 1923 1263 1957 1297
rect 483 1183 517 1217
rect 1923 1183 1957 1217
rect 1923 1103 1957 1137
rect 1343 943 1377 977
rect 2503 943 2537 977
rect 1193 753 1227 787
rect 1773 753 1807 787
rect 2503 523 2537 557
rect 2503 443 2537 477
rect 2503 363 2537 397
<< metal1 >>
rect 40 1900 2140 1980
rect 40 1490 120 1900
rect 900 1470 980 1900
rect 1480 1470 1560 1900
rect 2060 1490 2140 1900
rect 460 1297 540 1320
rect 460 1263 483 1297
rect 517 1280 540 1297
rect 1900 1297 1980 1320
rect 1900 1280 1923 1297
rect 517 1263 1923 1280
rect 1957 1263 1980 1297
rect 460 1240 1980 1263
rect 0 1160 390 1240
rect 460 1217 2880 1240
rect 460 1183 483 1217
rect 517 1200 1923 1217
rect 517 1183 540 1200
rect 460 1160 540 1183
rect 310 810 390 1160
rect 1170 787 1250 1200
rect 1900 1183 1923 1200
rect 1957 1183 2880 1217
rect 1900 1160 2880 1183
rect 1900 1137 1980 1160
rect 1900 1103 1923 1137
rect 1957 1103 1980 1137
rect 1900 1080 1980 1103
rect 1320 977 2560 1000
rect 1320 943 1343 977
rect 1377 943 2503 977
rect 2537 943 2560 977
rect 1320 920 2560 943
rect 1170 753 1193 787
rect 1227 753 1250 787
rect 1170 730 1250 753
rect 1750 787 1830 920
rect 1750 753 1773 787
rect 1807 753 1830 787
rect 1750 730 1830 753
rect 2330 500 2420 720
rect 0 420 2420 500
rect 2480 557 2560 580
rect 2480 523 2503 557
rect 2537 523 2560 557
rect 2480 500 2560 523
rect 2480 477 2880 500
rect 2480 443 2503 477
rect 2537 443 2880 477
rect 2480 420 2880 443
rect 2480 397 2560 420
rect 2480 363 2503 397
rect 2537 363 2560 397
rect 2480 340 2560 363
rect 40 -100 120 250
rect 900 -100 980 250
rect 1480 -100 1560 250
rect 2060 -100 2140 250
rect 40 -180 2140 -100
use dco_aux_inv  dco_aux_inv_0
timestamp 1729593089
transform 1 0 1120 0 1 880
box -260 -700 320 680
use dco_aux_inv  dco_aux_inv_1
timestamp 1729593089
transform 1 0 1700 0 1 880
box -260 -700 320 680
use dco_main_inv  dco_main_inv_0
timestamp 1729593089
transform 1 0 260 0 1 880
box -260 -880 600 860
use dco_main_inv  dco_main_inv_1
timestamp 1729593089
transform 1 0 2280 0 1 880
box -260 -880 600 860
<< labels >>
rlabel metal1 s 60 1980 60 1980 4 VCCA
rlabel locali s 1290 1740 1290 1740 4 VPWR
rlabel metal1 s 2880 1200 2880 1200 4 outp
rlabel metal1 s 0 1200 0 1200 4 inp
rlabel metal1 s 0 460 0 460 4 inn
rlabel metal1 s 2880 460 2880 460 4 outn
rlabel metal1 s 130 -180 130 -180 4 GND
rlabel locali s 1310 0 1310 0 4 VGND
<< end >>
