magic
tech sky130A
magscale 1 2
timestamp 1723886438
<< nwell >>
rect 3102 402 3218 722
rect 3102 400 3276 402
rect 1118 -400 1456 -78
rect 3645 -212 3825 -86
rect 3645 -214 3848 -212
rect 3645 -324 3836 -214
rect 3645 -332 3848 -324
rect 3645 -407 3825 -332
<< pwell >>
rect 3068 162 3280 298
rect 1094 -640 1494 -460
rect 3606 -494 3868 -466
rect 3604 -552 3868 -494
rect 3606 -646 3868 -552
rect 3608 -654 3866 -646
<< psubdiff >>
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 3140 188 3202 224
rect 1128 -526 1190 -494
rect 1128 -560 1144 -526
rect 1178 -560 1190 -526
rect 1128 -594 1190 -560
rect 3676 -596 3776 -582
rect 3676 -630 3712 -596
rect 3746 -630 3776 -596
rect 3676 -644 3776 -630
<< nsubdiff >>
rect 3136 564 3198 592
rect 3136 530 3148 564
rect 3182 530 3198 564
rect 3136 492 3198 530
rect 1156 -274 1218 -242
rect 1156 -308 1172 -274
rect 1206 -308 1218 -274
rect 1156 -342 1218 -308
rect 3780 -258 3836 -224
rect 3780 -292 3794 -258
rect 3828 -292 3836 -258
rect 3780 -324 3836 -292
<< psubdiffcont >>
rect 3156 224 3190 258
rect 1144 -560 1178 -526
rect 3712 -630 3746 -596
<< nsubdiffcont >>
rect 3148 530 3182 564
rect 1172 -308 1206 -274
rect 3794 -292 3828 -258
<< locali >>
rect 3136 564 3198 592
rect 3136 530 3148 564
rect 3182 530 3198 564
rect 3136 492 3198 530
rect 1446 352 1560 462
rect 2258 352 2380 462
rect 3072 352 3270 458
rect 3966 352 4084 462
rect 4776 352 4894 462
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 3140 188 3202 224
rect 1156 -274 1218 -242
rect 1156 -308 1172 -274
rect 1206 -308 1218 -274
rect 1156 -342 1218 -308
rect 3780 -258 3836 -224
rect 3780 -292 3794 -258
rect 3828 -292 3836 -258
rect 3780 -324 3836 -292
rect 1128 -526 1190 -494
rect 1128 -560 1144 -526
rect 1178 -560 1190 -526
rect 1128 -594 1190 -560
rect 3676 -596 3776 -582
rect 3676 -630 3712 -596
rect 3746 -630 3776 -596
rect 3676 -644 3776 -630
<< viali >>
rect 3148 530 3182 564
rect 5530 468 5564 502
rect 810 368 844 402
rect 3156 224 3190 258
rect 948 -286 982 -252
rect 1172 -308 1206 -274
rect 3794 -292 3828 -258
rect 1516 -444 1550 -410
rect 3368 -444 3402 -410
rect 3538 -454 3572 -420
rect 3900 -452 3934 -418
rect 3990 -456 4024 -422
rect 1768 -500 1802 -466
rect 1144 -560 1178 -526
rect 2880 -538 2914 -504
rect 3454 -562 3488 -528
rect 3712 -630 3746 -596
<< metal1 >>
rect 3136 564 3198 592
rect 3136 530 3148 564
rect 3182 530 3198 564
rect 3136 492 3198 530
rect 5514 540 5590 548
rect 5514 502 5948 540
rect 5514 468 5530 502
rect 5564 468 5948 502
rect 746 434 886 464
rect 5514 440 5948 468
rect 444 402 886 434
rect 444 374 810 402
rect 444 38 504 374
rect 746 368 810 374
rect 844 368 886 402
rect 746 350 886 368
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 3140 188 3202 224
rect 5848 58 5948 440
rect 444 -22 1402 38
rect 934 -252 994 -202
rect 934 -286 948 -252
rect 982 -286 994 -252
rect 934 -372 994 -286
rect 1156 -274 1218 -242
rect 1156 -308 1172 -274
rect 1206 -308 1218 -274
rect 1156 -342 1218 -308
rect 1342 -338 1402 -22
rect 3676 -42 5948 58
rect 936 -392 994 -372
rect 936 -452 1312 -392
rect 1342 -398 1572 -338
rect 1128 -526 1190 -494
rect 1128 -560 1144 -526
rect 1178 -560 1190 -526
rect 1128 -594 1190 -560
rect 1266 -510 1312 -452
rect 1502 -410 1572 -398
rect 3676 -402 3736 -42
rect 3780 -258 3836 -224
rect 3780 -292 3794 -258
rect 3828 -292 3836 -258
rect 3780 -324 3836 -292
rect 1502 -444 1516 -410
rect 1550 -444 1572 -410
rect 1502 -468 1572 -444
rect 3122 -410 3418 -402
rect 3122 -444 3368 -410
rect 3402 -444 3418 -410
rect 1758 -466 1814 -452
rect 1758 -500 1768 -466
rect 1802 -500 1814 -466
rect 3122 -458 3418 -444
rect 3518 -420 3736 -402
rect 3518 -454 3538 -420
rect 3572 -454 3736 -420
rect 3122 -496 3192 -458
rect 3518 -462 3736 -454
rect 3798 -418 3950 -402
rect 3798 -452 3900 -418
rect 3934 -452 3950 -418
rect 3518 -472 3576 -462
rect 3798 -470 3950 -452
rect 3984 -422 4212 -406
rect 3984 -456 3990 -422
rect 4024 -456 4212 -422
rect 3984 -468 4212 -456
rect 3798 -494 3858 -470
rect 1758 -510 1814 -500
rect 1266 -570 1814 -510
rect 2862 -504 3192 -496
rect 3604 -504 3858 -494
rect 2862 -538 2880 -504
rect 2914 -538 3192 -504
rect 2862 -570 3192 -538
rect 3444 -528 3858 -504
rect 3444 -562 3454 -528
rect 3488 -552 3858 -528
rect 3488 -562 3604 -552
rect 3444 -564 3604 -562
rect 3444 -580 3500 -564
rect 3676 -596 3776 -582
rect 3676 -630 3712 -596
rect 3746 -630 3776 -596
rect 3676 -644 3776 -630
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 730 0 1 -662
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1484 0 1 -662
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 730 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_1
timestamp 1701704242
transform 1 0 1542 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_2
timestamp 1701704242
transform 1 0 2354 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_3
timestamp 1701704242
transform 1 0 3248 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_4
timestamp 1701704242
transform 1 0 4060 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_5
timestamp 1701704242
transform 1 0 4872 0 1 140
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3862 0 1 -668
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3332 0 1 -668
box -38 -48 314 592
<< end >>
