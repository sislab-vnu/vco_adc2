magic
tech sky130A
timestamp 1725397606
<< nwell >>
rect -60 1080 2805 1105
rect -60 925 -40 1080
rect 0 1070 1935 1080
rect 0 1060 910 1070
rect 950 1060 1390 1070
rect 1430 1060 1935 1070
rect 0 925 895 1060
rect -60 885 895 925
rect 1695 925 1935 1060
rect 1975 970 2805 1080
rect 1975 925 2710 970
rect 1695 885 2710 925
rect -60 550 2710 885
rect -60 515 1795 550
rect -60 505 1670 515
rect 1835 505 2710 550
<< pwell >>
rect -60 470 1670 480
rect -60 440 1795 470
rect 1835 440 2710 480
rect -60 160 0 440
rect 815 160 2710 440
rect -60 -20 -40 160
rect 815 40 910 160
rect 0 0 910 40
rect 950 5 1390 160
rect 1430 5 1935 160
rect 1975 120 2710 160
rect 1975 5 2805 120
rect 950 0 2805 5
rect 0 -20 2805 0
<< psubdiff >>
rect 840 150 880 165
rect 840 130 850 150
rect 870 130 880 150
rect 840 110 880 130
rect 840 90 850 110
rect 870 90 880 110
rect 840 70 880 90
rect 840 50 850 70
rect 870 50 880 70
rect 840 35 880 50
rect 1865 150 1905 165
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 1865 110 1905 130
rect 1865 90 1875 110
rect 1895 90 1905 110
rect 1865 70 1905 90
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 1865 35 1905 50
<< nsubdiff >>
rect 840 1035 880 1050
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 840 995 880 1015
rect 840 975 850 995
rect 870 975 880 995
rect 840 955 880 975
rect 840 935 850 955
rect 870 935 880 955
rect 840 920 880 935
rect 1865 1045 1905 1060
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 1865 1005 1905 1025
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 1865 965 1905 985
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 1865 930 1905 945
<< psubdiffcont >>
rect 850 130 870 150
rect 850 90 870 110
rect 850 50 870 70
rect 1875 130 1895 150
rect 1875 90 1895 110
rect 1875 50 1895 70
<< nsubdiffcont >>
rect 850 1015 870 1035
rect 850 975 870 995
rect 850 935 870 955
rect 1875 1025 1895 1045
rect 1875 985 1895 1005
rect 1875 945 1895 965
<< polycont >>
rect 1090 480 1110 500
rect 1130 480 1150 500
rect 1170 480 1190 500
rect 1560 480 1580 500
rect 1600 480 1620 500
rect 1640 480 1660 500
<< locali >>
rect 735 1135 2040 1175
rect 840 1035 880 1135
rect 910 1050 950 1135
rect 1390 1050 1430 1135
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 840 995 880 1015
rect 840 975 850 995
rect 870 975 880 995
rect 840 955 880 975
rect 840 935 850 955
rect 870 935 880 955
rect 840 920 880 935
rect 1865 1045 1905 1135
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 1865 1005 1905 1025
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 1865 965 1905 985
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 1865 930 1905 945
rect 405 650 655 680
rect 625 505 655 650
rect 1080 505 1200 525
rect 1550 505 1670 525
rect 625 500 1200 505
rect 625 480 1090 500
rect 1110 480 1130 500
rect 1150 480 1170 500
rect 1190 480 1200 500
rect 625 475 1200 480
rect 1355 500 1670 505
rect 1355 480 1560 500
rect 1580 480 1600 500
rect 1620 480 1640 500
rect 1660 480 1670 500
rect 1355 475 1670 480
rect 1080 460 1200 475
rect 1550 460 1670 475
rect 840 150 880 165
rect 840 130 850 150
rect 870 130 880 150
rect 840 110 880 130
rect 840 90 850 110
rect 870 90 880 110
rect 840 70 880 90
rect 840 50 850 70
rect 870 50 880 70
rect 840 35 880 50
rect 1865 150 1905 165
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 1865 110 1905 130
rect 1865 90 1875 110
rect 1895 90 1905 110
rect 1865 70 1905 90
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 910 -50 950 40
rect 1390 -50 1430 40
rect 1865 35 1905 50
rect 575 -90 1970 -50
<< viali >>
rect 850 1015 870 1035
rect 850 975 870 995
rect 850 935 870 955
rect 1875 1025 1895 1045
rect 1875 985 1895 1005
rect 1875 945 1895 965
rect 375 775 395 795
rect 1805 780 1825 800
rect 1090 480 1110 500
rect 1130 480 1150 500
rect 1170 480 1190 500
rect 1560 480 1580 500
rect 1600 480 1620 500
rect 1640 480 1660 500
rect 1325 250 1345 270
rect 2350 250 2370 270
rect 850 130 870 150
rect 850 90 870 110
rect 850 50 870 70
rect 1875 130 1895 150
rect 1875 90 1895 110
rect 1875 50 1895 70
<< metal1 >>
rect 840 1035 880 1125
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 840 995 880 1015
rect 840 975 850 995
rect 870 975 880 995
rect 840 955 880 975
rect 840 935 850 955
rect 870 935 880 955
rect 840 920 880 935
rect 1865 1045 1905 1125
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 1865 1005 1905 1025
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 1865 965 1905 985
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 1865 930 1905 945
rect -60 765 190 815
rect 365 800 2805 815
rect 365 795 1805 800
rect 365 775 375 795
rect 395 780 1805 795
rect 1825 780 2805 800
rect 395 775 2805 780
rect 365 765 2805 775
rect 140 525 190 765
rect 835 615 2105 665
rect 835 290 885 615
rect 2055 525 2105 615
rect 1080 500 1200 525
rect 1080 480 1090 500
rect 1110 480 1130 500
rect 1150 480 1170 500
rect 1190 480 1200 500
rect 1080 460 1200 480
rect 1550 500 1670 525
rect 1550 480 1560 500
rect 1580 480 1600 500
rect 1620 480 1640 500
rect 1660 480 1670 500
rect 1550 460 1670 480
rect 1585 290 1635 460
rect -60 240 885 290
rect 1315 270 2805 290
rect 1315 250 1325 270
rect 1345 250 2350 270
rect 2370 250 2805 270
rect 1315 240 2805 250
rect 840 150 880 165
rect 840 130 850 150
rect 870 130 880 150
rect 840 120 880 130
rect 1865 150 1905 165
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 1865 120 1905 130
rect 840 110 1905 120
rect 840 90 850 110
rect 870 90 1875 110
rect 1895 90 1905 110
rect 840 80 1905 90
rect 840 70 880 80
rect 840 50 850 70
rect 870 50 880 70
rect 840 -40 880 50
rect 1865 70 1905 80
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 1865 -40 1905 50
use aux_inv_vco  aux_inv_vco_0
timestamp 1725396630
transform 1 0 885 0 1 500
box 0 -500 490 590
use aux_inv_vco  aux_inv_vco_1
timestamp 1725396630
transform 1 0 1365 0 1 500
box 0 -500 490 590
use main_inv_vco  main_inv_vco_0
timestamp 1725081791
transform 1 0 -1060 0 1 545
box 1000 -635 1890 630
use main_inv_vco  main_inv_vco_1
timestamp 1725081791
transform 1 0 915 0 1 545
box 1000 -635 1890 630
<< labels >>
rlabel metal1 2805 785 2805 785 3 OUT_P
port 3 e
rlabel metal1 2805 265 2805 265 3 OUT_N
port 4 e
rlabel locali 1410 1175 1410 1175 1 VPWR
port 5 n
rlabel locali 1410 -90 1410 -90 5 VGND
port 6 s
<< end >>
