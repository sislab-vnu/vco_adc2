* this file contains all digital circuits written by SPICE
