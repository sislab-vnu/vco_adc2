magic
tech sky130A
timestamp 1723605105
<< checkpaint >>
rect -630 -630 640 640
<< nwell >>
rect 0 0 10 10
<< pdiff >>
rect 2 2 8 8
<< end >>
