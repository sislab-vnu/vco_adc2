** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/cc_inv.sch
.subckt cc_inv inp inn outp outn VGND VDDA GND
*.PININFO outp:O inn:I VGND:B outn:O inp:I VDDA:B GND:B
Xi_1 inp outp VGND VDDA GND main_inv
Xi_2 inn outn VGND VDDA GND main_inv
Xi_3 outp outn VGND VDDA GND aux_inv
Xi_4 outn outp VGND VDDA GND aux_inv
.ends

* expanding   symbol:  main_inv.sym # of pins=5
** sym_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sym
** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sch
.subckt main_inv A Y VGND VDDA GND
*.PININFO VDDA:B VGND:B A:I Y:O GND:B
XM2 Y A VGND GND sky130_fd_pr__nfet_01v8 L=3.65 W=8 nf=2 m=1
XM1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=10 nf=2 m=1
.ends


* expanding   symbol:  aux_inv.sym # of pins=5
** sym_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sym
** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sch
.subckt aux_inv A Y VGND VDDA GND
*.PININFO VDDA:B VGND:B A:I Y:O GND:B
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=3.65 W=4 nf=1 m=1
XM2 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=5 nf=1 m=1
.ends

.end
