* NGSPICE file created from ring_osc.ext - technology: sky130A

.subckt main_inv_vco a_0_n1090# a_1540_n1010# a_730_0# a_n80_n1010# a_1540_0# w_n120_n40#
+ a_n80_0# VSUBS
X0 a_1540_0# a_0_n1090# a_730_0# w_n120_n40# sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65
X1 a_730_n1010# a_0_n1090# a_n80_n1010# VSUBS sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65
X2 a_1540_n1010# a_0_n1090# a_730_n1010# VSUBS sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=3.65
X3 a_730_0# a_0_n1090# a_n80_0# w_n120_n40# sky130_fd_pr__pfet_01v8 ad=1 pd=5.4 as=2 ps=10.8 w=5 l=3.65
.ends

.subckt inv a_0_n1090# a_730_0# a_n80_n1010# w_n120_n40# a_730_n1010# a_n80_0# VSUBS
X0 a_730_n1010# a_0_n1090# a_n80_n1010# VSUBS sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
X1 a_730_0# a_0_n1090# a_n80_0# w_n120_n40# sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
.ends

.subckt cc_inv inp inn outp GND VPWR VGND VCCA
Xmain_inv_vco_1 inn outp li_4680_1990# VGND outp VCCA VPWR GND main_inv_vco
Xmain_inv_vco_0 inp outp main_inv_vco_0/a_730_0# VGND outp VCCA VPWR GND main_inv_vco
Xinv_2 outp outp VGND VCCA outp VPWR GND inv
Xinv_3 outp outp VGND VCCA outp VPWR GND inv
.ends

.subckt ring_osc
Xcc_inv_0 cc_inv_0/inp cc_inv_0/inp cc_inv_1/inp VSUBS cc_inv_0/VPWR VSUBS cc_inv_2/VCCA
+ cc_inv
Xcc_inv_2 cc_inv_2/inp cc_inv_2/inp cc_inv_4/inp VSUBS cc_inv_2/VPWR VSUBS cc_inv_2/VCCA
+ cc_inv
Xcc_inv_1 cc_inv_1/inp cc_inv_1/inp cc_inv_2/inp VSUBS cc_inv_1/VPWR VSUBS cc_inv_2/VCCA
+ cc_inv
Xcc_inv_3 cc_inv_3/inp cc_inv_3/inp cc_inv_0/inp VSUBS cc_inv_3/VPWR VSUBS cc_inv_4/VCCA
+ cc_inv
Xcc_inv_4 cc_inv_4/inp cc_inv_4/inp cc_inv_3/inp VSUBS cc_inv_4/VPWR VSUBS cc_inv_4/VCCA
+ cc_inv
.ends

