magic
tech sky130A
timestamp 1723696154
<< pwell >>
rect -60 -20 290 200
<< nmos >>
rect 0 0 50 180
rect 90 0 140 180
rect 180 0 230 180
<< ndiff >>
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 90 90 110
rect 50 70 60 90
rect 80 70 90 90
rect 50 50 90 70
rect 50 30 60 50
rect 80 30 90 50
rect 50 0 90 30
rect 140 170 180 180
rect 140 150 150 170
rect 170 150 180 170
rect 140 130 180 150
rect 140 110 150 130
rect 170 110 180 130
rect 140 90 180 110
rect 140 70 150 90
rect 170 70 180 90
rect 140 50 180 70
rect 140 30 150 50
rect 170 30 180 50
rect 140 0 180 30
rect 230 170 270 180
rect 230 150 240 170
rect 260 150 270 170
rect 230 130 270 150
rect 230 110 240 130
rect 260 110 270 130
rect 230 90 270 110
rect 230 70 240 90
rect 260 70 270 90
rect 230 50 270 70
rect 230 30 240 50
rect 260 30 270 50
rect 230 0 270 30
<< ndiffc >>
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 60 150 80 170
rect 60 110 80 130
rect 60 70 80 90
rect 60 30 80 50
rect 150 150 170 170
rect 150 110 170 130
rect 150 70 170 90
rect 150 30 170 50
rect 240 150 260 170
rect 240 110 260 130
rect 240 70 260 90
rect 240 30 260 50
<< poly >>
rect 0 180 50 200
rect 90 180 140 200
rect 180 180 230 200
rect 0 -20 50 0
rect 90 -20 140 0
rect 180 -20 230 0
<< locali >>
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 90 90 110
rect 50 70 60 90
rect 80 70 90 90
rect 50 50 90 70
rect 50 30 60 50
rect 80 30 90 50
rect 50 0 90 30
rect 140 170 180 180
rect 140 150 150 170
rect 170 150 180 170
rect 140 130 180 150
rect 140 110 150 130
rect 170 110 180 130
rect 140 90 180 110
rect 140 70 150 90
rect 170 70 180 90
rect 140 50 180 70
rect 140 30 150 50
rect 170 30 180 50
rect 140 0 180 30
rect 230 170 270 180
rect 230 150 240 170
rect 260 150 270 170
rect 230 130 270 150
rect 230 110 240 130
rect 260 110 270 130
rect 230 90 270 110
rect 230 70 240 90
rect 260 70 270 90
rect 230 50 270 70
rect 230 30 240 50
rect 260 30 270 50
rect 230 0 270 30
<< end >>
