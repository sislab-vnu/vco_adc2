* NGSPICE file created from DLib_UpDownCounter.ext - technology: sky130A





.subckt DLib_UpDownCounter UP DOWN setB Dout_buf VDDA GND
Xsky130_fd_sc_hd__dfstp_1_0 UP_buf Q2N SetBi GND GND VDDA VDDA Q1 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfstp_1_1 DWN_buf Q1_buf SetBi GND GND VDDA VDDA Q2 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__inv_2_0 setB GND GND VDDA VDDA SetBi sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_1 DOWN GND GND VDDA VDDA DWN_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_1 Q2 GND GND VDDA VDDA Q2N sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_2 Dout GND GND VDDA VDDA Dout_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_3 Q1 GND GND VDDA VDDA Q1_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_4 UP GND GND VDDA VDDA UP_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_1 Q1 Q2 GND GND VDDA VDDA Dout sky130_fd_sc_hd__xor2_1
.ends


