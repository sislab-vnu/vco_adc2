* NGSPICE file created from dco_idac.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_R469US a_n35_840# VSUBS
X0 a_n35_840# a_n35_n1272# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

*.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
*.subckt sky130_fd_sc_hd__buf_2 1   2   3   4   5   6
.subckt sky130_fd_sc_hd__buf_2 1 2 3 4 5 6
X0 5 a_27_47# 6 4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR 1 a_27_47# 4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 6 a_27_47# 2 3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15 M=2
X3 2 1 a_27_47# 3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

*.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
*.subckt sky130_fd_sc_hd__inv_2 1  2    3   4   5   6
.subckt sky130_fd_sc_hd__inv_2 1 2 3 4 5 6
X0 6 1 5 4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15 M=2
X1 2 1 6 3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
.ends

.subckt dco_idac Dctrl Vbs1 Vbs2 Vbs3 Vbs4 Isup
Xsky130_fd_pr__res_xhigh_po_0p35_R469US_0 Isup Isup sky130_fd_pr__res_xhigh_po_0p35_R469US
Xsky130_fd_sc_hd__buf_2_0 Dctrl sky130_fd_sc_hd__buf_2_0/VGND Isup sky130_fd_sc_hd__buf_2_0/VPB
+ sky130_fd_sc_hd__buf_2_0/VPWR sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/VGND
+ Isup sky130_fd_sc_hd__inv_2_0/VPB sky130_fd_sc_hd__inv_2_0/VPWR sky130_fd_sc_hd__inv_2_0/Y
+ sky130_fd_sc_hd__inv_2
X0 w_n580_n1630# sky130_fd_sc_hd__inv_2_0/A Isup w_n580_n1630# sky130_fd_pr__pfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.5 M=2
X1 Isup sky130_fd_sc_hd__inv_2_0/A w_n580_n1630# Isup sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X2 w_2370_n90# Vbs1 w_n580_n80# w_n580_n80# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X3 w_n580_n1630# Vbs4 w_1270_n80# w_1270_n80# sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X4 Isup sky130_fd_sc_hd__inv_2_0/Y w_n580_n1630# Isup sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X5 w_1270_n80# Vbs3 w_n580_n80# w_n580_n80# sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X6 Isup Vbs2 w_2370_n90# w_2370_n90# sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X7 Isup sky130_fd_sc_hd__inv_2_0/Y w_n580_n1630# w_n580_n1630# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
.ends

