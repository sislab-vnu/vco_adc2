magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -260 -90 850 1070
<< pwell >>
rect -106 -904 836 -194
rect -246 -1046 836 -904
rect -246 -1056 -114 -1046
<< nmos >>
rect 0 -1020 730 -220
<< pmos >>
rect 0 -10 730 990
<< ndiff >>
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -643 0 -597
rect -80 -677 -57 -643
rect -23 -677 0 -643
rect -80 -723 0 -677
rect -80 -757 -57 -723
rect -23 -757 0 -723
rect -80 -803 0 -757
rect -80 -837 -57 -803
rect -23 -837 0 -803
rect -80 -883 0 -837
rect -80 -917 -57 -883
rect -23 -917 0 -883
rect -80 -963 0 -917
rect -80 -997 -57 -963
rect -23 -997 0 -963
rect -80 -1020 0 -997
rect 730 -243 810 -220
rect 730 -277 753 -243
rect 787 -277 810 -243
rect 730 -323 810 -277
rect 730 -357 753 -323
rect 787 -357 810 -323
rect 730 -403 810 -357
rect 730 -437 753 -403
rect 787 -437 810 -403
rect 730 -483 810 -437
rect 730 -517 753 -483
rect 787 -517 810 -483
rect 730 -563 810 -517
rect 730 -597 753 -563
rect 787 -597 810 -563
rect 730 -643 810 -597
rect 730 -677 753 -643
rect 787 -677 810 -643
rect 730 -723 810 -677
rect 730 -757 753 -723
rect 787 -757 810 -723
rect 730 -803 810 -757
rect 730 -837 753 -803
rect 787 -837 810 -803
rect 730 -883 810 -837
rect 730 -917 753 -883
rect 787 -917 810 -883
rect 730 -963 810 -917
rect 730 -997 753 -963
rect 787 -997 810 -963
rect 730 -1020 810 -997
<< pdiff >>
rect -80 967 0 990
rect -80 933 -57 967
rect -23 933 0 967
rect -80 887 0 933
rect -80 853 -57 887
rect -23 853 0 887
rect -80 807 0 853
rect -80 773 -57 807
rect -23 773 0 807
rect -80 727 0 773
rect -80 693 -57 727
rect -23 693 0 727
rect -80 647 0 693
rect -80 613 -57 647
rect -23 613 0 647
rect -80 567 0 613
rect -80 533 -57 567
rect -23 533 0 567
rect -80 487 0 533
rect -80 453 -57 487
rect -23 453 0 487
rect -80 407 0 453
rect -80 373 -57 407
rect -23 373 0 407
rect -80 327 0 373
rect -80 293 -57 327
rect -23 293 0 327
rect -80 247 0 293
rect -80 213 -57 247
rect -23 213 0 247
rect -80 167 0 213
rect -80 133 -57 167
rect -23 133 0 167
rect -80 87 0 133
rect -80 53 -57 87
rect -23 53 0 87
rect -80 -10 0 53
rect 730 967 810 990
rect 730 933 753 967
rect 787 933 810 967
rect 730 887 810 933
rect 730 853 753 887
rect 787 853 810 887
rect 730 807 810 853
rect 730 773 753 807
rect 787 773 810 807
rect 730 727 810 773
rect 730 693 753 727
rect 787 693 810 727
rect 730 647 810 693
rect 730 613 753 647
rect 787 613 810 647
rect 730 567 810 613
rect 730 533 753 567
rect 787 533 810 567
rect 730 487 810 533
rect 730 453 753 487
rect 787 453 810 487
rect 730 407 810 453
rect 730 373 753 407
rect 787 373 810 407
rect 730 327 810 373
rect 730 293 753 327
rect 787 293 810 327
rect 730 247 810 293
rect 730 213 753 247
rect 787 213 810 247
rect 730 167 810 213
rect 730 133 753 167
rect 787 133 810 167
rect 730 87 810 133
rect 730 53 753 87
rect 787 53 810 87
rect 730 -10 810 53
<< ndiffc >>
rect -57 -277 -23 -243
rect -57 -357 -23 -323
rect -57 -437 -23 -403
rect -57 -517 -23 -483
rect -57 -597 -23 -563
rect -57 -677 -23 -643
rect -57 -757 -23 -723
rect -57 -837 -23 -803
rect -57 -917 -23 -883
rect -57 -997 -23 -963
rect 753 -277 787 -243
rect 753 -357 787 -323
rect 753 -437 787 -403
rect 753 -517 787 -483
rect 753 -597 787 -563
rect 753 -677 787 -643
rect 753 -757 787 -723
rect 753 -837 787 -803
rect 753 -917 787 -883
rect 753 -997 787 -963
<< pdiffc >>
rect -57 933 -23 967
rect -57 853 -23 887
rect -57 773 -23 807
rect -57 693 -23 727
rect -57 613 -23 647
rect -57 533 -23 567
rect -57 453 -23 487
rect -57 373 -23 407
rect -57 293 -23 327
rect -57 213 -23 247
rect -57 133 -23 167
rect -57 53 -23 87
rect 753 933 787 967
rect 753 853 787 887
rect 753 773 787 807
rect 753 693 787 727
rect 753 613 787 647
rect 753 533 787 567
rect 753 453 787 487
rect 753 373 787 407
rect 753 293 787 327
rect 753 213 787 247
rect 753 133 787 167
rect 753 53 787 87
<< psubdiff >>
rect -220 -963 -140 -930
rect -220 -997 -197 -963
rect -163 -997 -140 -963
rect -220 -1030 -140 -997
<< nsubdiff >>
rect -220 967 -140 1000
rect -220 933 -197 967
rect -163 933 -140 967
rect -220 900 -140 933
<< psubdiffcont >>
rect -197 -997 -163 -963
<< nsubdiffcont >>
rect -197 933 -163 967
<< poly >>
rect 0 990 730 1070
rect 0 -220 730 -10
rect 0 -1100 730 -1020
<< locali >>
rect -220 967 -140 1000
rect -220 933 -197 967
rect -163 933 -140 967
rect -220 900 -140 933
rect -80 967 0 990
rect -80 933 -57 967
rect -23 933 0 967
rect -80 887 0 933
rect -80 853 -57 887
rect -23 853 0 887
rect -80 807 0 853
rect -80 773 -57 807
rect -23 773 0 807
rect -80 727 0 773
rect -80 693 -57 727
rect -23 693 0 727
rect -80 647 0 693
rect -80 613 -57 647
rect -23 613 0 647
rect -80 567 0 613
rect -80 533 -57 567
rect -23 533 0 567
rect -80 487 0 533
rect -80 453 -57 487
rect -23 453 0 487
rect -80 407 0 453
rect -80 373 -57 407
rect -23 373 0 407
rect -80 327 0 373
rect -80 293 -57 327
rect -23 293 0 327
rect -80 247 0 293
rect -80 213 -57 247
rect -23 213 0 247
rect -80 167 0 213
rect -80 133 -57 167
rect -23 133 0 167
rect -80 87 0 133
rect -80 53 -57 87
rect -23 53 0 87
rect -80 -10 0 53
rect 730 967 810 990
rect 730 933 753 967
rect 787 933 810 967
rect 730 887 810 933
rect 730 853 753 887
rect 787 853 810 887
rect 730 807 810 853
rect 730 773 753 807
rect 787 773 810 807
rect 730 727 810 773
rect 730 693 753 727
rect 787 693 810 727
rect 730 647 810 693
rect 730 613 753 647
rect 787 613 810 647
rect 730 567 810 613
rect 730 533 753 567
rect 787 533 810 567
rect 730 487 810 533
rect 730 453 753 487
rect 787 453 810 487
rect 730 407 810 453
rect 730 373 753 407
rect 787 373 810 407
rect 730 327 810 373
rect 730 293 753 327
rect 787 293 810 327
rect 730 247 810 293
rect 730 213 753 247
rect 787 213 810 247
rect 730 167 810 213
rect 730 133 753 167
rect 787 133 810 167
rect 730 87 810 133
rect 730 53 753 87
rect 787 53 810 87
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -643 0 -597
rect -80 -677 -57 -643
rect -23 -677 0 -643
rect -80 -723 0 -677
rect -80 -757 -57 -723
rect -23 -757 0 -723
rect -80 -803 0 -757
rect -80 -837 -57 -803
rect -23 -837 0 -803
rect -80 -883 0 -837
rect -80 -917 -57 -883
rect -23 -917 0 -883
rect -220 -963 -140 -930
rect -220 -997 -197 -963
rect -163 -997 -140 -963
rect -220 -1030 -140 -997
rect -80 -963 0 -917
rect -80 -997 -57 -963
rect -23 -997 0 -963
rect -80 -1020 0 -997
rect 730 -243 810 53
rect 730 -277 753 -243
rect 787 -277 810 -243
rect 730 -323 810 -277
rect 730 -357 753 -323
rect 787 -357 810 -323
rect 730 -403 810 -357
rect 730 -437 753 -403
rect 787 -437 810 -403
rect 730 -483 810 -437
rect 730 -517 753 -483
rect 787 -517 810 -483
rect 730 -563 810 -517
rect 730 -597 753 -563
rect 787 -597 810 -563
rect 730 -643 810 -597
rect 730 -677 753 -643
rect 787 -677 810 -643
rect 730 -723 810 -677
rect 730 -757 753 -723
rect 787 -757 810 -723
rect 730 -803 810 -757
rect 730 -837 753 -803
rect 787 -837 810 -803
rect 730 -883 810 -837
rect 730 -917 753 -883
rect 787 -917 810 -883
rect 730 -963 810 -917
rect 730 -997 753 -963
rect 787 -997 810 -963
rect 730 -1020 810 -997
<< viali >>
rect -197 933 -163 967
rect -197 -997 -163 -963
<< metal1 >>
rect -220 967 -140 1000
rect -220 933 -197 967
rect -163 933 -140 967
rect -220 900 -140 933
rect -220 -963 -140 -930
rect -220 -997 -197 -963
rect -163 -997 -140 -963
rect -220 -1030 -140 -997
<< labels >>
rlabel poly s 0 -120 0 -120 4 A
rlabel locali s -40 990 -40 990 4 VPWR
rlabel locali s -40 -1020 -40 -1020 4 VGND
rlabel locali s 810 -120 810 -120 4 Y
rlabel metal1 s -180 1000 -180 1000 4 VCCA
rlabel metal1 s -180 -1030 -180 -1030 4 GND
<< end >>
