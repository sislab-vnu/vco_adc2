magic
tech sky130A
timestamp 1723711581
<< nwell >>
rect -60 -20 110 200
<< pmos >>
rect 0 0 50 180
<< pdiff >>
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 90 90 110
rect 50 70 60 90
rect 80 70 90 90
rect 50 50 90 70
rect 50 30 60 50
rect 80 30 90 50
rect 50 0 90 30
<< pdiffc >>
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 60 150 80 170
rect 60 110 80 130
rect 60 70 80 90
rect 60 30 80 50
<< poly >>
rect 0 180 50 200
rect 0 -20 50 0
<< locali >>
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 90 90 110
rect 50 70 60 90
rect 80 70 90 90
rect 50 50 90 70
rect 50 30 60 50
rect 80 30 90 50
rect 50 0 90 30
<< end >>
