magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect 3080 3500 3256 3820
rect 7210 900 7340 1220
<< pwell >>
rect 3152 3250 3266 3402
rect 7204 674 7316 826
<< psubdiff >>
rect 3178 3342 3240 3376
rect 3178 3308 3195 3342
rect 3229 3308 3240 3342
rect 3178 3276 3240 3308
rect 7230 767 7290 800
rect 7230 733 7243 767
rect 7277 733 7290 767
rect 7230 700 7290 733
<< nsubdiff >>
rect 3160 3662 3220 3696
rect 3160 3628 3174 3662
rect 3208 3628 3220 3662
rect 3160 3596 3220 3628
rect 7230 1017 7290 1050
rect 7230 983 7243 1017
rect 7277 983 7290 1017
rect 7230 950 7290 983
<< psubdiffcont >>
rect 3195 3308 3229 3342
rect 7243 733 7277 767
<< nsubdiffcont >>
rect 3174 3628 3208 3662
rect 7243 983 7277 1017
<< locali >>
rect 2600 5897 2640 5900
rect 2600 5863 2603 5897
rect 2637 5863 2640 5897
rect 2600 5860 2640 5863
rect 3180 5897 3220 5900
rect 3180 5863 3183 5897
rect 3217 5863 3220 5897
rect 3180 5860 3220 5863
rect 3760 5897 3800 5900
rect 3760 5863 3763 5897
rect 3797 5863 3800 5897
rect 3760 5860 3800 5863
rect 4620 5897 4660 5900
rect 4620 5863 4623 5897
rect 4657 5863 4660 5897
rect 4620 5860 4660 5863
rect 5480 5897 5520 5900
rect 5480 5863 5483 5897
rect 5517 5863 5520 5897
rect 5480 5860 5520 5863
rect 6060 5897 6100 5900
rect 6060 5863 6063 5897
rect 6097 5863 6100 5897
rect 6060 5860 6100 5863
rect 6640 5897 6680 5900
rect 6640 5863 6643 5897
rect 6677 5863 6680 5897
rect 6640 5860 6680 5863
rect 7500 5897 7540 5900
rect 7500 5863 7503 5897
rect 7537 5863 7540 5897
rect 7500 5860 7540 5863
rect 8360 5897 8400 5900
rect 8360 5863 8363 5897
rect 8397 5863 8400 5897
rect 8360 5860 8400 5863
rect 8940 5897 8980 5900
rect 8940 5863 8943 5897
rect 8977 5863 8980 5897
rect 8940 5860 8980 5863
rect 9520 5897 9560 5900
rect 9520 5863 9523 5897
rect 9557 5863 9560 5897
rect 9520 5860 9560 5863
rect 2600 4237 2640 4240
rect 2600 4203 2603 4237
rect 2637 4203 2640 4237
rect 2600 4200 2640 4203
rect 3180 4237 3220 4240
rect 3180 4203 3183 4237
rect 3217 4203 3220 4237
rect 3180 4200 3220 4203
rect 3760 4237 3800 4240
rect 3760 4203 3763 4237
rect 3797 4203 3800 4237
rect 3760 4200 3800 4203
rect 4620 4237 4660 4240
rect 4620 4203 4623 4237
rect 4657 4203 4660 4237
rect 4620 4200 4660 4203
rect 5480 4237 5520 4240
rect 5480 4203 5483 4237
rect 5517 4203 5520 4237
rect 5480 4200 5520 4203
rect 6060 4237 6100 4240
rect 6060 4203 6063 4237
rect 6097 4203 6100 4237
rect 6060 4200 6100 4203
rect 6640 4237 6680 4240
rect 6640 4203 6643 4237
rect 6677 4203 6680 4237
rect 6640 4200 6680 4203
rect 7500 4237 7540 4240
rect 7500 4203 7503 4237
rect 7537 4203 7540 4237
rect 7500 4200 7540 4203
rect 8360 4237 8400 4240
rect 8360 4203 8363 4237
rect 8397 4203 8400 4237
rect 8360 4200 8400 4203
rect 8940 4237 8980 4240
rect 8940 4203 8943 4237
rect 8977 4203 8980 4237
rect 8940 4200 8980 4203
rect 3160 3667 3220 3696
rect 3730 3670 4190 3730
rect 3160 3633 3173 3667
rect 3207 3662 3220 3667
rect 3160 3628 3174 3633
rect 3208 3628 3220 3662
rect 3160 3596 3220 3628
rect 3330 3497 3370 3500
rect 3330 3463 3333 3497
rect 3367 3463 3370 3497
rect 3330 3460 3370 3463
rect 3690 3487 3760 3500
rect 3690 3453 3703 3487
rect 3737 3453 3760 3487
rect 3690 3440 3760 3453
rect 3170 3342 3240 3380
rect 3170 3308 3195 3342
rect 3229 3308 3240 3342
rect 3170 3170 3240 3308
rect 3290 3170 3360 3230
rect 3170 3100 3360 3170
rect 3170 2730 3270 3100
rect 4130 3040 4190 3670
rect 4400 3437 5390 3460
rect 4400 3403 5333 3437
rect 5367 3403 5390 3437
rect 4400 3380 5390 3403
rect 5910 3437 5950 3440
rect 5910 3403 5913 3437
rect 5947 3403 5950 3437
rect 5910 3400 5950 3403
rect 6490 3437 6530 3440
rect 6490 3403 6493 3437
rect 6527 3403 6530 3437
rect 6490 3400 6530 3403
rect 7350 3437 7390 3440
rect 7350 3403 7353 3437
rect 7387 3403 7390 3437
rect 7350 3400 7390 3403
rect 8210 3437 8250 3440
rect 8210 3403 8213 3437
rect 8247 3403 8250 3437
rect 8210 3400 8250 3403
rect 8790 3437 8830 3440
rect 8790 3403 8793 3437
rect 8827 3403 8830 3437
rect 8790 3400 8830 3403
rect 9370 3437 9410 3440
rect 9370 3403 9373 3437
rect 9407 3403 9410 3437
rect 9370 3400 9410 3403
rect 4120 3017 4200 3040
rect 4120 2983 4143 3017
rect 4177 2983 4200 3017
rect 4120 2960 4200 2983
rect 4400 2730 4480 3380
rect 3170 2650 4480 2730
rect 3170 1012 3270 2650
rect 5330 1777 5370 1780
rect 5330 1743 5333 1777
rect 5367 1743 5370 1777
rect 5330 1740 5370 1743
rect 5910 1777 5950 1780
rect 5910 1743 5913 1777
rect 5947 1743 5950 1777
rect 5910 1740 5950 1743
rect 6490 1777 6530 1780
rect 6490 1743 6493 1777
rect 6527 1743 6530 1777
rect 6490 1740 6530 1743
rect 7350 1777 7390 1780
rect 7350 1743 7353 1777
rect 7387 1743 7390 1777
rect 7350 1740 7390 1743
rect 8210 1777 8250 1780
rect 8210 1743 8213 1777
rect 8247 1743 8250 1777
rect 8210 1740 8250 1743
rect 8790 1777 8830 1780
rect 8790 1743 8793 1777
rect 8827 1743 8830 1777
rect 8790 1740 8830 1743
rect 9370 1777 9410 1780
rect 9370 1743 9373 1777
rect 9407 1743 9410 1777
rect 9370 1740 9410 1743
rect 10230 1777 10270 1780
rect 10230 1743 10233 1777
rect 10267 1743 10270 1777
rect 10230 1740 10270 1743
rect 3170 978 3198 1012
rect 3232 978 3270 1012
rect 3170 940 3270 978
rect 5980 1537 6080 1560
rect 5980 1503 6013 1537
rect 6047 1503 6080 1537
rect 2320 600 2510 680
rect 5980 -270 6080 1503
rect 7950 1357 8460 1390
rect 7950 1323 7983 1357
rect 8017 1323 8063 1357
rect 8097 1323 8143 1357
rect 8177 1323 8223 1357
rect 8257 1323 8303 1357
rect 8337 1323 8383 1357
rect 8417 1323 8460 1357
rect 7950 1290 8460 1323
rect 7230 1017 7290 1050
rect 7230 983 7243 1017
rect 7277 983 7290 1017
rect 7230 950 7290 983
rect 7230 767 7290 800
rect 7230 733 7243 767
rect 7277 733 7290 767
rect 7090 490 7170 630
rect 7230 490 7290 733
rect 7090 430 7290 490
rect 7950 480 8050 1290
rect 8360 630 8460 1290
rect 7090 250 7170 430
rect 7090 150 7620 250
rect 7090 110 7190 150
rect 8410 110 8440 120
rect 7090 30 8440 110
rect 7090 -2090 7190 30
rect 7090 -2190 7620 -2090
rect 7090 -2230 7190 -2190
rect 8410 -2230 8450 -2220
rect 7090 -2300 8450 -2230
rect 2750 -4080 2950 -3120
rect 7090 -4080 7190 -2300
rect 2750 -4280 7190 -4080
<< viali >>
rect 2603 5863 2637 5897
rect 3183 5863 3217 5897
rect 3763 5863 3797 5897
rect 4623 5863 4657 5897
rect 5483 5863 5517 5897
rect 6063 5863 6097 5897
rect 6643 5863 6677 5897
rect 7503 5863 7537 5897
rect 8363 5863 8397 5897
rect 8943 5863 8977 5897
rect 9523 5863 9557 5897
rect 2603 4203 2637 4237
rect 3183 4203 3217 4237
rect 3763 4203 3797 4237
rect 4623 4203 4657 4237
rect 5483 4203 5517 4237
rect 6063 4203 6097 4237
rect 6643 4203 6677 4237
rect 7503 4203 7537 4237
rect 8363 4203 8397 4237
rect 8943 4203 8977 4237
rect 3173 3662 3207 3667
rect 3173 3633 3174 3662
rect 3174 3633 3207 3662
rect 3333 3463 3367 3497
rect 3703 3453 3737 3487
rect 3195 3308 3229 3342
rect 5333 3403 5367 3437
rect 5913 3403 5947 3437
rect 6493 3403 6527 3437
rect 7353 3403 7387 3437
rect 8213 3403 8247 3437
rect 8793 3403 8827 3437
rect 9373 3403 9407 3437
rect 4143 2983 4177 3017
rect 5333 1743 5367 1777
rect 5913 1743 5947 1777
rect 6493 1743 6527 1777
rect 7353 1743 7387 1777
rect 8213 1743 8247 1777
rect 8793 1743 8827 1777
rect 9373 1743 9407 1777
rect 10233 1743 10267 1777
rect 3198 978 3232 1012
rect 6013 1503 6047 1537
rect 7983 1323 8017 1357
rect 8063 1323 8097 1357
rect 8143 1323 8177 1357
rect 8223 1323 8257 1357
rect 8303 1323 8337 1357
rect 8383 1323 8417 1357
rect 7028 1050 7062 1084
rect 7028 974 7062 1008
rect 7243 983 7277 1017
rect 6846 854 6880 888
rect 7243 733 7277 767
<< metal1 >>
rect 2600 5897 2640 5900
rect 2600 5863 2603 5897
rect 2637 5863 2640 5897
rect 2600 5860 2640 5863
rect 3180 5897 3220 5900
rect 3180 5863 3183 5897
rect 3217 5863 3220 5897
rect 3180 5860 3220 5863
rect 3760 5897 3800 5900
rect 3760 5863 3763 5897
rect 3797 5863 3800 5897
rect 3760 5860 3800 5863
rect 4620 5897 4660 5900
rect 4620 5863 4623 5897
rect 4657 5863 4660 5897
rect 4620 5860 4660 5863
rect 5480 5897 5520 5900
rect 5480 5863 5483 5897
rect 5517 5863 5520 5897
rect 5480 5860 5520 5863
rect 6060 5897 6100 5900
rect 6060 5863 6063 5897
rect 6097 5863 6100 5897
rect 6060 5860 6100 5863
rect 6640 5897 6680 5900
rect 6640 5863 6643 5897
rect 6677 5863 6680 5897
rect 6640 5860 6680 5863
rect 7500 5897 7540 5900
rect 7500 5863 7503 5897
rect 7537 5863 7540 5897
rect 7500 5860 7540 5863
rect 8360 5897 8400 5900
rect 8360 5863 8363 5897
rect 8397 5863 8400 5897
rect 8360 5860 8400 5863
rect 8940 5897 8980 5900
rect 8940 5863 8943 5897
rect 8977 5863 8980 5897
rect 8940 5860 8980 5863
rect 9520 5897 9560 5900
rect 9520 5863 9523 5897
rect 9557 5863 9560 5897
rect 9520 5860 9560 5863
rect 4520 5340 4740 5420
rect 2600 4237 2640 4240
rect 2600 4203 2603 4237
rect 2637 4203 2640 4237
rect 2600 4200 2640 4203
rect 3180 4237 3220 4240
rect 3180 4203 3183 4237
rect 3217 4203 3220 4237
rect 3180 4200 3220 4203
rect 3760 4237 3800 4240
rect 3760 4203 3763 4237
rect 3797 4203 3800 4237
rect 3760 4200 3800 4203
rect 4620 4237 4660 4240
rect 4620 4203 4623 4237
rect 4657 4203 4660 4237
rect 4620 4200 4660 4203
rect 5480 4237 5520 4240
rect 5480 4203 5483 4237
rect 5517 4203 5520 4237
rect 5480 4200 5520 4203
rect 6060 4237 6100 4240
rect 6060 4203 6063 4237
rect 6097 4203 6100 4237
rect 6060 4200 6100 4203
rect 6640 4237 6680 4240
rect 6640 4203 6643 4237
rect 6677 4203 6680 4237
rect 6640 4200 6680 4203
rect 7500 4237 7540 4240
rect 7500 4203 7503 4237
rect 7537 4203 7540 4237
rect 7500 4200 7540 4203
rect 8360 4237 8400 4240
rect 8360 4203 8363 4237
rect 8397 4203 8400 4237
rect 8360 4200 8400 4203
rect 8940 4237 8980 4240
rect 8940 4203 8943 4237
rect 8977 4203 8980 4237
rect 8940 4200 8980 4203
rect 3160 3816 3300 3830
rect 3160 3764 3174 3816
rect 3226 3764 3300 3816
rect 3160 3740 3300 3764
rect 3920 3806 4010 3830
rect 3920 3754 3944 3806
rect 3996 3754 4010 3806
rect 3160 3667 3220 3740
rect 3160 3633 3173 3667
rect 3207 3633 3220 3667
rect 3160 3596 3220 3633
rect 3300 3497 3400 3540
rect 3920 3500 4010 3754
rect 3300 3490 3333 3497
rect 2890 3463 3333 3490
rect 3367 3463 3400 3497
rect 2890 3430 3400 3463
rect 3680 3487 4010 3500
rect 3680 3453 3703 3487
rect 3737 3453 4010 3487
rect 3680 3430 4010 3453
rect 5330 3437 5370 3440
rect 5330 3403 5333 3437
rect 5367 3403 5370 3437
rect 5330 3400 5370 3403
rect 5910 3437 5950 3440
rect 5910 3403 5913 3437
rect 5947 3403 5950 3437
rect 5910 3400 5950 3403
rect 6490 3437 6530 3440
rect 6490 3403 6493 3437
rect 6527 3403 6530 3437
rect 6490 3400 6530 3403
rect 7350 3437 7390 3440
rect 7350 3403 7353 3437
rect 7387 3403 7390 3437
rect 7350 3400 7390 3403
rect 8210 3437 8250 3440
rect 8210 3403 8213 3437
rect 8247 3403 8250 3437
rect 8210 3400 8250 3403
rect 8790 3437 8830 3440
rect 8790 3403 8793 3437
rect 8827 3403 8830 3437
rect 8790 3400 8830 3403
rect 9370 3437 9410 3440
rect 9370 3403 9373 3437
rect 9407 3403 9410 3437
rect 9370 3400 9410 3403
rect 3178 3342 3240 3376
rect 3178 3308 3195 3342
rect 3229 3308 3240 3342
rect 3178 3276 3240 3308
rect 4140 3017 4180 3020
rect 4140 2983 4143 3017
rect 4177 2983 4180 3017
rect 4140 2980 4180 2983
rect 4220 1240 4300 2280
rect 5330 1777 5370 1780
rect 5330 1743 5333 1777
rect 5367 1743 5370 1777
rect 5330 1740 5370 1743
rect 5910 1777 5950 1780
rect 5910 1743 5913 1777
rect 5947 1743 5950 1777
rect 5910 1740 5950 1743
rect 6490 1777 6530 1780
rect 6490 1743 6493 1777
rect 6527 1743 6530 1777
rect 6490 1740 6530 1743
rect 7350 1777 7390 1780
rect 7350 1743 7353 1777
rect 7387 1743 7390 1777
rect 7350 1740 7390 1743
rect 8210 1777 8250 1780
rect 8210 1743 8213 1777
rect 8247 1743 8250 1777
rect 8210 1740 8250 1743
rect 8790 1777 8830 1780
rect 8790 1743 8793 1777
rect 8827 1743 8830 1777
rect 8790 1740 8830 1743
rect 9370 1777 9410 1780
rect 9370 1743 9373 1777
rect 9407 1743 9410 1777
rect 9370 1740 9410 1743
rect 10230 1777 10270 1780
rect 10230 1743 10233 1777
rect 10267 1743 10270 1777
rect 10230 1740 10270 1743
rect 6010 1537 6050 1540
rect 6010 1503 6013 1537
rect 6047 1503 6050 1537
rect 6010 1500 6050 1503
rect 7180 1376 7290 1390
rect 7180 1324 7214 1376
rect 7266 1324 7290 1376
rect 4220 1160 6490 1240
rect 7180 1230 7290 1324
rect 7950 1366 8460 1390
rect 7950 1314 7974 1366
rect 8026 1357 8134 1366
rect 8186 1357 8294 1366
rect 8346 1357 8460 1366
rect 8026 1323 8063 1357
rect 8097 1323 8134 1357
rect 8186 1323 8223 1357
rect 8257 1323 8294 1357
rect 8346 1323 8383 1357
rect 8417 1323 8460 1357
rect 8026 1314 8134 1323
rect 8186 1314 8294 1323
rect 8346 1314 8460 1323
rect 7950 1290 8460 1314
rect 3170 1012 6270 1040
rect 3170 978 3198 1012
rect 3232 978 6270 1012
rect 3170 940 6270 978
rect 2540 770 5590 870
rect 2540 480 2640 770
rect 3960 480 4060 590
rect 3750 380 4390 480
rect 5490 470 5590 770
rect 6170 250 6270 940
rect 6410 910 6490 1160
rect 7160 1140 7290 1230
rect 7020 1084 7070 1100
rect 7020 1050 7028 1084
rect 7062 1050 7070 1084
rect 7020 1008 7070 1050
rect 7020 974 7028 1008
rect 7062 974 7070 1008
rect 6410 908 6830 910
rect 6410 888 6896 908
rect 6410 854 6846 888
rect 6880 854 6896 888
rect 7020 900 7070 974
rect 7230 1017 7290 1140
rect 7230 983 7243 1017
rect 7277 983 7290 1017
rect 7230 950 7290 983
rect 7350 900 8270 930
rect 7020 860 8270 900
rect 7037 858 8270 860
rect 6410 836 6896 854
rect 6410 830 6830 836
rect 7350 830 8270 858
rect 7230 767 7290 800
rect 7230 733 7243 767
rect 7277 733 7290 767
rect 7230 700 7290 733
rect 8170 350 8270 830
rect 6170 150 7540 250
rect 11080 -74 11180 -50
rect 11080 -126 11104 -74
rect 11156 -126 11180 -74
rect 11080 -150 11180 -126
rect 11840 -74 11940 -50
rect 11840 -126 11864 -74
rect 11916 -126 11940 -74
rect 1240 -1540 1320 -1340
rect 1540 -1364 1640 -1340
rect 1540 -1416 1564 -1364
rect 1616 -1416 1640 -1364
rect 1540 -1480 1640 -1416
rect 11840 -1430 11940 -126
rect 8140 -1530 11940 -1430
rect 6530 -1784 7730 -1760
rect 6530 -1836 6554 -1784
rect 6606 -1836 7730 -1784
rect 6530 -1860 7730 -1836
rect 8040 -1860 8050 -1760
rect 8140 -1960 8240 -1530
rect 11080 -2414 11180 -2390
rect 11080 -2466 11104 -2414
rect 11156 -2466 11180 -2414
rect 7680 -2580 7930 -2490
rect 11080 -2500 11180 -2466
<< via1 >>
rect 3174 3764 3226 3816
rect 3944 3754 3996 3806
rect 7214 1324 7266 1376
rect 7974 1357 8026 1366
rect 8134 1357 8186 1366
rect 8294 1357 8346 1366
rect 7974 1323 7983 1357
rect 7983 1323 8017 1357
rect 8017 1323 8026 1357
rect 8134 1323 8143 1357
rect 8143 1323 8177 1357
rect 8177 1323 8186 1357
rect 8294 1323 8303 1357
rect 8303 1323 8337 1357
rect 8337 1323 8346 1357
rect 7974 1314 8026 1323
rect 8134 1314 8186 1323
rect 8294 1314 8346 1323
rect 11104 -126 11156 -74
rect 11864 -126 11916 -74
rect 1564 -1416 1616 -1364
rect 6554 -1836 6606 -1784
rect 11104 -2466 11156 -2414
<< metal2 >>
rect 3130 3816 4010 3830
rect 3130 3764 3174 3816
rect 3226 3806 4010 3816
rect 3226 3764 3944 3806
rect 3130 3754 3944 3764
rect 3996 3754 4010 3806
rect 3130 3740 4010 3754
rect 3920 1390 4010 3740
rect 1540 1376 8460 1390
rect 1540 1324 7214 1376
rect 7266 1366 8460 1376
rect 7266 1324 7974 1366
rect 1540 1314 7974 1324
rect 8026 1314 8134 1366
rect 8186 1314 8294 1366
rect 8346 1314 8460 1366
rect 1540 1300 8460 1314
rect 1540 -1364 1640 1300
rect 1540 -1416 1564 -1364
rect 1616 -1416 1640 -1364
rect 1540 -1440 1640 -1416
rect 6530 -1784 6630 1300
rect 7950 1290 8460 1300
rect 11080 -74 11940 -50
rect 11080 -126 11104 -74
rect 11156 -126 11864 -74
rect 11916 -126 11940 -74
rect 11080 -150 11940 -126
rect 6530 -1836 6554 -1784
rect 6606 -1836 6630 -1784
rect 6530 -1860 6630 -1836
rect 11080 -2414 11890 -2390
rect 11080 -2466 11104 -2414
rect 11156 -2466 11890 -2414
rect 11080 -2490 11890 -2466
use dco_freq  dco_freq_0
timestamp 1729593089
transform 1 0 8320 0 1 50
box -880 -1250 3330 640
use dco_freq  dco_freq_1
timestamp 1729593089
transform 1 0 8320 0 1 -2290
box -880 -1250 3330 640
use dco_idac  dco_idac_0
timestamp 1729593089
transform 1 0 2860 0 1 -60
box -1860 -3150 3220 740
use dco_ring_osc  dco_ring_osc_0
timestamp 1729593089
transform 1 0 1680 0 1 4000
box -500 -2520 9440 2160
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0
timestamp 1729593089
transform 1 0 6808 0 1 638
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0
timestamp 1729593089
transform 1 0 3288 0 1 3238
box -38 -48 498 592
<< labels >>
rlabel locali s 6040 1560 6040 1560 4 Isup
rlabel metal2 s 11900 -50 11900 -50 4 ro_div2
rlabel metal1 s 7560 930 7560 930 4 pha_ro
rlabel metal1 s 4340 1240 4340 1240 4 p_osc
rlabel metal2 s 1580 1390 1580 1390 4 VCCD
rlabel locali s 2380 680 2380 680 4 VCCA
rlabel metal1 s 1290 -1340 1290 -1340 4 Dctrl
rlabel metal1 s 2930 3490 2930 3490 4 ENB
rlabel metal1 s 2700 870 2700 870 4 Vbs_12
rlabel metal1 s 4010 590 4010 590 4 Vbs_34
rlabel metal2 s 11820 -2390 11820 -2390 4 pha_DCO
rlabel locali s 4910 -4080 4910 -4080 4 GND
<< end >>
