magic
tech sky130A
timestamp 1726043895
<< nwell >>
rect -130 -40 160 340
<< pwell >>
rect -130 -350 160 -70
<< nmos >>
rect 0 -310 100 -110
<< pmos >>
rect 0 0 100 300
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -310 0 -300
rect 100 -120 140 -110
rect 100 -140 110 -120
rect 130 -140 140 -120
rect 100 -160 140 -140
rect 100 -180 110 -160
rect 130 -180 140 -160
rect 100 -200 140 -180
rect 100 -220 110 -200
rect 130 -220 140 -200
rect 100 -240 140 -220
rect 100 -260 110 -240
rect 130 -260 140 -240
rect 100 -280 140 -260
rect 100 -300 110 -280
rect 130 -300 140 -280
rect 100 -310 140 -300
<< pdiff >>
rect -40 290 0 300
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 100 290 140 300
rect 100 270 110 290
rect 130 270 140 290
rect 100 250 140 270
rect 100 230 110 250
rect 130 230 140 250
rect 100 210 140 230
rect 100 190 110 210
rect 130 190 140 210
rect 100 170 140 190
rect 100 150 110 170
rect 130 150 140 170
rect 100 130 140 150
rect 100 110 110 130
rect 130 110 140 130
rect 100 90 140 110
rect 100 70 110 90
rect 130 70 140 90
rect 100 50 140 70
rect 100 30 110 50
rect 130 30 140 50
rect 100 0 140 30
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect 110 -140 130 -120
rect 110 -180 130 -160
rect 110 -220 130 -200
rect 110 -260 130 -240
rect 110 -300 130 -280
<< pdiffc >>
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 110 270 130 290
rect 110 230 130 250
rect 110 190 130 210
rect 110 150 130 170
rect 110 110 130 130
rect 110 70 130 90
rect 110 30 130 50
<< psubdiff >>
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< nsubdiff >>
rect -110 280 -70 295
rect -110 260 -100 280
rect -80 260 -70 280
rect -110 245 -70 260
<< psubdiffcont >>
rect -100 -300 -80 -280
<< nsubdiffcont >>
rect -100 260 -80 280
<< poly >>
rect 0 300 100 340
rect 0 -110 100 0
rect 0 -350 100 -310
<< locali >>
rect -110 280 -70 295
rect -110 260 -100 280
rect -80 260 -70 280
rect -110 245 -70 260
rect -40 290 0 300
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 100 290 140 300
rect 100 270 110 290
rect 130 270 140 290
rect 100 250 140 270
rect 100 230 110 250
rect 130 230 140 250
rect 100 210 140 230
rect 100 190 110 210
rect 130 190 140 210
rect 100 170 140 190
rect 100 150 110 170
rect 130 150 140 170
rect 100 130 140 150
rect 100 110 110 130
rect 130 110 140 130
rect 100 90 140 110
rect 100 70 110 90
rect 130 70 140 90
rect 100 50 140 70
rect 100 30 110 50
rect 130 30 140 50
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -310 0 -300
rect 100 -120 140 30
rect 100 -140 110 -120
rect 130 -140 140 -120
rect 100 -160 140 -140
rect 100 -180 110 -160
rect 130 -180 140 -160
rect 100 -200 140 -180
rect 100 -220 110 -200
rect 130 -220 140 -200
rect 100 -240 140 -220
rect 100 -260 110 -240
rect 130 -260 140 -240
rect 100 -280 140 -260
rect 100 -300 110 -280
rect 130 -300 140 -280
rect 100 -310 140 -300
<< viali >>
rect -100 260 -80 280
rect -100 -300 -80 -280
<< metal1 >>
rect -110 280 -70 295
rect -110 260 -100 280
rect -80 260 -70 280
rect -110 245 -70 260
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< labels >>
rlabel locali -20 300 -20 300 1 VPWR
port 1 n
rlabel metal1 -90 295 -90 295 1 VCCA
port 2 n
rlabel poly 0 -55 0 -55 7 A
port 3 w
rlabel locali 140 -55 140 -55 3 Y
port 4 e
rlabel metal1 -90 -265 -90 -265 1 GND
port 5 n
rlabel locali -20 -310 -20 -310 5 VGND
port 6 s
<< end >>
