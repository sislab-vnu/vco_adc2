magic
tech sky130A
magscale 1 2
timestamp 1727170671
<< locali >>
rect -2760 4470 2150 4580
rect -2740 4170 -2480 4270
rect -2740 4100 -2650 4170
rect -2580 4150 -2480 4170
rect -2580 4110 3220 4150
rect -2580 4100 3130 4110
rect -2740 4070 3130 4100
rect 3170 4070 3220 4110
rect -2740 4050 3220 4070
rect -2740 4010 -2480 4050
rect -4470 3590 2990 3650
rect -4470 -1750 -4410 3590
rect -4470 -1830 1430 -1750
rect -4470 -3890 -4410 -1830
rect -3300 -2860 -3200 -2830
rect -3300 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3300 -2920 -3200 -2900
rect 1350 -3350 1430 -1830
rect 15700 -1800 15770 -1070
rect 15700 -1840 15720 -1800
rect 15760 -1840 15770 -1800
rect 15700 -1860 15770 -1840
rect 19560 -2490 21710 -2480
rect 19560 -2530 19580 -2490
rect 19620 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 19560 -2550 21710 -2530
rect 18400 -3200 18470 -2660
rect 1350 -3370 5570 -3350
rect 1350 -3410 5520 -3370
rect 5560 -3410 5570 -3370
rect 1350 -3430 5570 -3410
rect -4470 -3930 -4460 -3890
rect -4420 -3930 -4410 -3890
rect -4470 -11680 -4410 -3930
rect 390 -4850 570 -4820
rect 390 -4890 500 -4850
rect 540 -4890 570 -4850
rect 390 -4920 570 -4890
rect 2700 -6190 4920 -6170
rect 2700 -6230 2720 -6190
rect 2760 -6230 4920 -6190
rect 2700 -6250 4920 -6230
rect 14840 -7240 15030 -7200
rect 14840 -7270 15490 -7240
rect 14840 -7320 14910 -7270
rect 14960 -7320 15490 -7270
rect 14840 -7380 15030 -7320
rect 15280 -8300 15380 -8270
rect 15280 -8340 15310 -8300
rect 15350 -8340 15380 -8300
rect 9710 -11000 10040 -10930
rect 9710 -11060 9740 -11000
rect 9800 -11060 9920 -11000
rect 9980 -11060 10040 -11000
rect 9710 -11130 10040 -11060
rect 15280 -11680 15380 -8340
rect 19080 -9260 19180 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 19180 -9260
rect 19080 -9330 19180 -9300
rect -4470 -11780 15380 -11680
<< viali >>
rect 540 7650 580 7690
rect 1630 7650 1670 7690
rect 2720 7650 2760 7690
rect 4640 7650 4680 7690
rect 6540 7650 6580 7690
rect 7630 7650 7670 7690
rect 8720 7650 8760 7690
rect 10640 7650 10680 7690
rect 12540 7650 12580 7690
rect 13630 7650 13670 7690
rect 14720 7650 14760 7690
rect 17420 7650 17460 7690
rect -2650 4100 -2580 4170
rect 3130 4070 3170 4110
rect 6400 1000 6440 1040
rect 7490 1000 7530 1040
rect 8580 1000 8620 1040
rect 10480 1000 10520 1040
rect 12400 1000 12440 1040
rect 13490 1000 13530 1040
rect 14580 1000 14620 1040
rect 16480 1000 16520 1040
rect 17420 1000 17460 1040
rect 740 -2610 780 -2570
rect -3270 -2900 -3230 -2860
rect 15720 -1840 15760 -1800
rect 19580 -2530 19620 -2490
rect 21650 -2530 21690 -2490
rect 5520 -3410 5560 -3370
rect -4460 -3930 -4420 -3890
rect 500 -4890 540 -4850
rect 2720 -6230 2760 -6190
rect 14910 -7320 14960 -7270
rect 15310 -8340 15350 -8300
rect 9740 -11060 9800 -11000
rect 9920 -11060 9980 -11000
rect 19110 -9300 19150 -9260
<< metal1 >>
rect -2080 7910 -1310 8010
rect -2740 4200 -2480 4270
rect -2740 4070 -2680 4200
rect -2550 4070 -2480 4200
rect -2740 4010 -2480 4070
rect -3390 1560 -1760 1660
rect -3390 -2830 -3300 1560
rect 6380 -60 6460 890
rect 13640 680 13740 710
rect 2700 -140 6460 -60
rect 730 -2560 1240 -2550
rect 730 -2570 780 -2560
rect 730 -2610 740 -2570
rect 730 -2620 780 -2610
rect 840 -2620 1240 -2560
rect 730 -2630 1240 -2620
rect -3390 -2860 -3200 -2830
rect -3390 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3390 -2920 -3200 -2900
rect -3390 -3056 -3280 -3050
rect -3390 -3080 -3060 -3056
rect -3390 -3140 -3370 -3080
rect -3310 -3140 -3060 -3080
rect -3390 -3156 -3060 -3140
rect -3390 -3160 -3280 -3156
rect -4470 -3890 -3160 -3870
rect -4470 -3930 -4460 -3890
rect -4420 -3930 -3160 -3890
rect -4470 -3950 -3160 -3930
rect -70 -3970 60 -3960
rect -70 -4030 -10 -3970
rect 50 -4030 60 -3970
rect -70 -4040 60 -4030
rect 470 -4850 570 -4820
rect 470 -4890 500 -4850
rect 540 -4890 570 -4850
rect 470 -12490 570 -4890
rect 2700 -6190 2780 -140
rect 6380 -720 6460 -690
rect 13640 -1070 13740 -690
rect 14930 -1600 15640 -1500
rect 5500 -3370 5570 -3350
rect 5500 -3410 5520 -3370
rect 5560 -3410 5570 -3370
rect 5500 -3430 5570 -3410
rect 14930 -5475 15030 -1600
rect 19560 -2490 19640 -2470
rect 19560 -2530 19580 -2490
rect 19620 -2530 19640 -2490
rect 19560 -2550 19640 -2530
rect 21610 -2490 21710 -2480
rect 21610 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 15480 -2640 15800 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2690 15800 -2640
rect 15560 -2700 15580 -2690
rect 15480 -2720 15580 -2700
rect 19930 -2860 20070 -2820
rect 19930 -2920 19970 -2860
rect 20030 -2920 20070 -2860
rect 19930 -2960 20070 -2920
rect 10995 -5565 15720 -5475
rect 3130 -5900 5260 -5800
rect 5160 -5960 5260 -5900
rect 2700 -6230 2720 -6190
rect 2760 -6230 2780 -6190
rect 2700 -6250 2780 -6230
rect 6580 -6300 6680 -6190
rect 15630 -6940 15720 -5565
rect 14840 -7260 15030 -7200
rect 14840 -7330 14900 -7260
rect 14970 -7330 15030 -7260
rect 14840 -7380 15030 -7330
rect 15280 -8286 15380 -8270
rect 15280 -8300 15570 -8286
rect 15280 -8340 15310 -8300
rect 15350 -8340 15570 -8300
rect 15280 -8356 15570 -8340
rect 15280 -8370 15380 -8356
rect 18700 -8376 18800 -8360
rect 18540 -8380 18800 -8376
rect 18540 -8440 18720 -8380
rect 18780 -8440 18800 -8380
rect 18540 -8446 18800 -8440
rect 18700 -8460 18800 -8446
rect 15830 -8920 15930 -8900
rect 15830 -8980 15850 -8920
rect 15910 -8980 15930 -8920
rect 15830 -9000 15930 -8980
rect 21610 -9230 21710 -2530
rect 19080 -9260 21710 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 21710 -9260
rect 19080 -9330 21710 -9300
rect 3420 -9970 3550 -9950
rect 3420 -9980 3630 -9970
rect 3420 -10040 3450 -9980
rect 3510 -10040 3630 -9980
rect 3420 -10050 3630 -10040
rect 3420 -10080 3550 -10050
rect 9710 -10980 10040 -10930
rect 9710 -11000 9820 -10980
rect 9710 -11060 9740 -11000
rect 9800 -11060 9820 -11000
rect 9710 -11070 9820 -11060
rect 9910 -11000 10040 -10980
rect 9910 -11060 9920 -11000
rect 9980 -11060 10040 -11000
rect 9910 -11070 10040 -11060
rect 9710 -11130 10040 -11070
rect 21610 -12490 21710 -9330
rect 470 -12590 21710 -12490
<< via1 >>
rect -1360 4900 -1300 4960
rect -2680 4170 -2550 4200
rect -2680 4100 -2650 4170
rect -2650 4100 -2580 4170
rect -2580 4100 -2550 4170
rect -2680 4070 -2550 4100
rect 780 -2620 840 -2560
rect -3370 -3140 -3310 -3080
rect -10 -4030 50 -3970
rect 15500 -2700 15560 -2640
rect 19970 -2920 20030 -2860
rect 14900 -7270 14970 -7260
rect 14900 -7320 14910 -7270
rect 14910 -7320 14960 -7270
rect 14960 -7320 14970 -7270
rect 14900 -7330 14970 -7320
rect 3870 -8260 3930 -8200
rect 18720 -8440 18780 -8380
rect 15850 -8980 15910 -8920
rect 3450 -10040 3510 -9980
rect 9820 -11070 9910 -10980
<< metal2 >>
rect -4970 4960 -1280 4980
rect -4970 4900 -1360 4960
rect -1300 4900 -1280 4960
rect -4970 4880 -1280 4900
rect -4970 -3050 -4870 4880
rect -2740 4200 -2480 4270
rect -2740 4070 -2680 4200
rect -2550 4070 -2480 4200
rect -2740 4010 -2480 4070
rect -2705 -165 -2515 4010
rect -2705 -355 2090 -165
rect 1900 -1085 2090 -355
rect 730 -2560 2000 -2550
rect 730 -2620 780 -2560
rect 840 -2620 2000 -2560
rect 730 -2630 2000 -2620
rect 15480 -2640 15580 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2700 15580 -2640
rect -5285 -3080 -3280 -3050
rect -5285 -3140 -3370 -3080
rect -3310 -3140 -3280 -3080
rect -5285 -3160 -3280 -3140
rect -4970 -9950 -4870 -3160
rect -20 -3970 1000 -3960
rect -20 -4030 -10 -3970
rect 50 -4030 1000 -3970
rect -20 -4040 1000 -4030
rect 920 -7670 1000 -4040
rect 15480 -6300 15580 -2700
rect 19930 -2860 20070 -2820
rect 19930 -2920 19970 -2860
rect 20030 -2920 20070 -2860
rect 19930 -2960 20070 -2920
rect 15480 -6400 19700 -6300
rect 14840 -7260 15030 -7200
rect 14840 -7330 14900 -7260
rect 14970 -7330 15030 -7260
rect 14840 -7380 15030 -7330
rect 920 -7750 3940 -7670
rect 3860 -8180 3940 -7750
rect 3850 -8200 3950 -8180
rect 3850 -8260 3870 -8200
rect 3930 -8260 3950 -8200
rect 3850 -8270 3950 -8260
rect 14869 -9240 14972 -7380
rect 19600 -8360 19700 -6400
rect 18700 -8380 19700 -8360
rect 18700 -8440 18720 -8380
rect 18780 -8440 19700 -8380
rect 18700 -8460 19700 -8440
rect 14330 -9340 14972 -9240
rect 14869 -9341 14972 -9340
rect 15120 -8900 15930 -8800
rect -4970 -9980 3550 -9950
rect -4970 -10040 3450 -9980
rect 3510 -10040 3550 -9980
rect -4970 -10080 3550 -10040
rect 9710 -10980 10040 -10930
rect 9710 -11070 9820 -10980
rect 9910 -11000 10040 -10980
rect 15120 -11000 15220 -8900
rect 15830 -8920 15930 -8900
rect 15830 -8980 15850 -8920
rect 15910 -8980 15930 -8920
rect 15830 -9000 15930 -8980
rect 19930 -11000 20030 -2960
rect 9910 -11070 20030 -11000
rect 9710 -11100 20030 -11070
rect 9710 -11130 10040 -11100
use count  count_0 ./../count
timestamp 1727161985
transform 1 0 -2340 0 1 -2076
box -880 -3154 3140 -440
use count  count_1
timestamp 1727161985
transform 1 0 16330 0 1 -6486
box -880 -3154 3140 -440
use dco  dco_0 ./../dco
timestamp 1727163546
transform 1 0 2620 0 1 -6850
box -720 -4280 11940 6160
use qz  qz_0 ./../quantizer
timestamp 1727164310
transform 1 0 15260 0 1 -2230
box 190 -710 5890 730
use vco  vco_0 ./../vco
timestamp 1727146712
transform 1 0 -2020 0 1 680
box 0 0 19930 7330
<< labels >>
rlabel metal1 6380 160 6380 160 7 VCCA
port 8 w
rlabel locali -2630 4580 -2630 4580 1 Anlg_in
port 3 n
rlabel metal2 -2620 4270 -2620 4270 1 VCCD
port 4 n
rlabel locali -3160 3650 -3160 3650 1 ENB
port 5 n
rlabel locali 15740 -1070 15740 -1070 1 CLK
port 2 n
rlabel locali 18400 -3160 18400 -3160 7 Dout
port 1 w
rlabel metal1 3300 -5800 3300 -5800 1 Vbs_12
port 7 n
rlabel metal1 6630 -6190 6630 -6190 1 Vbs_34
port 9 n
rlabel metal2 -5180 -3050 -5180 -3050 1 GND
port 6 n
rlabel metal2 3480 -7670 3480 -7670 1 D1
rlabel metal2 14720 -9240 14720 -9240 1 p_dco
<< end >>
