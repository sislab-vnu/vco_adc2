* NGSPICE file created from ALib_IDAC.ext - technology: sky130A



.subckt sky130_fd_pr__res_xhigh_po_0p35_RSCMUS a_n35_n1272# a_n35_840# a_n165_n1402#
X0 a_n35_840# a_n35_n1272# a_n165_n1402# sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

.subckt ALib_IDAC Vbs1 Vbs2 Vbs3 Vbs4 Dctrl Isup VDDA GND
Xsky130_fd_sc_hd__buf_2_0 Dctrl GND GND VDDA VDDA sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A GND GND VDDA VDDA sky130_fd_sc_hd__inv_2_0/Y
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0 GND a_n150_n1850# GND sky130_fd_pr__res_xhigh_po_0p35_RSCMUS
X0 Isup sky130_fd_sc_hd__inv_2_0/A w_n510_n1930# GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X1 w_2370_n90# Vbs1 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X2 w_n510_n1930# Vbs4 w_1270_n80# w_1270_n80# sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X3 a_n150_n1850# sky130_fd_sc_hd__inv_2_0/Y w_n510_n1930# GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X4 Isup sky130_fd_sc_hd__inv_2_0/Y w_n510_n1930# w_n510_n1930# sky130_fd_pr__pfet_01v8_hvt ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
X5 w_1270_n80# Vbs3 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X6 Isup Vbs2 w_2370_n90# w_2370_n90# sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X7 w_n510_n1930# sky130_fd_sc_hd__inv_2_0/A a_n150_n1850# w_n510_n1930# sky130_fd_pr__pfet_01v8_hvt ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.5 M=2
.ends


