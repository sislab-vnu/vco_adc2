* NGSPICE file created from idac.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_R469US a_n35_n1272# a_n35_840# VSUBS
X0 a_n35_840# a_n35_n1272# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

*.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
*.subckt sky130_fd_sc_hd__buf_2 1   2   3   4   5   6
.subckt sky130_fd_sc_hd__buf_2 1 2 3 4 5 6
X0 5 a_27_47# 6 4 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR 1 a_27_47# 4 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 6 a_27_47# 2 3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15 M=2
X3 2 1 a_27_47# 3 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

*.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
*.subckt sky130_fd_sc_hd__inv_2 1  2    3   4   5   6
.subckt sky130_fd_sc_hd__inv_2 1 2 3 4 5 6
X0 6 1 5 4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15 M=2
X1 2 1 6 3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
.ends

.subckt n_lk G S D B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5 M=2
.ends

.subckt p_lk G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
.ends

.subckt ol1 add_pwr g1 g2 VSUBS
Xn_lk_0 g2 VSUBS add_pwr VSUBS n_lk
Xp_lk_0 g1 add_pwr VSUBS add_pwr p_lk
.ends

.subckt p_br1 G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
.ends

.subckt p_br2 G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
.ends

.subckt obr s_1 g_1 d_1 s_2 g_2 d_2
Xp_br1_0 g_1 s_1 d_1 s_1 p_br1
Xp_br2_0 g_2 s_2 d_2 s_2 p_br2
.ends

.subckt idac
Xsky130_fd_pr__res_xhigh_po_0p35_R469US_0 obr_1/d_1 obr_1/d_1 obr_1/d_1 sky130_fd_pr__res_xhigh_po_0p35_R469US
Xsky130_fd_sc_hd__inv_2_0 ol1_1/g2 obr_1/d_1 obr_1/d_1 sky130_fd_sc_hd__inv_2_0/VPB
+ sky130_fd_sc_hd__inv_2_0/VPB ol1_1/g1 sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_0 sky130_fd_sc_hd__buf_2_0/A obr_1/d_1 obr_1/d_1 sky130_fd_sc_hd__inv_2_0/VPB
+ sky130_fd_sc_hd__inv_2_0/VPB ol1_1/g2 sky130_fd_sc_hd__buf_2
Xol1_0 obr_1/d_2 ol1_1/g2 ol1_1/g1 obr_1/d_1 ol1
Xol1_1 obr_1/d_2 ol1_1/g1 ol1_1/g2 obr_1/d_1 ol1
Xobr_1 obr_1/s_1 obr_1/g_1 obr_1/d_1 obr_1/s_2 obr_1/g_2 obr_1/d_2 obr
Xobr_0 obr_0/s_2 obr_0/g_1 obr_1/s_1 obr_0/s_2 obr_0/g_2 obr_1/s_2 obr
.ends

