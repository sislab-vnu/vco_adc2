magic
tech sky130A
magscale 1 2
timestamp 1723567583
<< pwell >>
rect 2590 1330 3100 1620
<< poly >>
rect 2000 2690 2080 2710
rect 2000 2650 2020 2690
rect 2060 2650 2080 2690
rect 2000 2500 2080 2650
rect 1790 2430 2080 2500
rect 2000 2330 2080 2430
rect 1790 2260 2080 2330
<< polycont >>
rect 2020 2650 2060 2690
<< viali >>
rect 2020 2650 2060 2690
rect 2663 1123 2697 1157
<< metal1 >>
rect 2000 2690 2080 2710
rect 2000 2650 2020 2690
rect 2060 2650 2080 2690
rect 2000 2630 2080 2650
rect 2454 1175 2554 1699
rect 2454 1157 2728 1175
rect 2454 1123 2663 1157
rect 2697 1123 2728 1157
rect 2454 1111 2728 1123
use ring_osc  ring_osc_0
timestamp 1723549246
transform 1 0 200 0 1 3020
box -340 -3020 17350 2290
use sky130_fd_pr__res_generic_po_C4R5Y4  sky130_fd_pr__res_generic_po_C4R5Y4_0
timestamp 1723566019
transform 0 1 1195 -1 0 2293
box -33 -595 33 595
use sky130_fd_pr__res_generic_po_C4R5Y4  sky130_fd_pr__res_generic_po_C4R5Y4_1
timestamp 1723566019
transform 0 1 1195 -1 0 2463
box -33 -595 33 595
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 3088 0 -1 1532
box -38 -48 498 592
<< end >>
