magic
tech sky130A
magscale 1 2
timestamp 1726807257
<< nwell >>
rect 7210 900 7340 1220
rect -410 -1130 -234 -810
<< pwell >>
rect 7170 660 7340 840
rect -334 -1372 -200 -1236
<< psubdiff >>
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7230 700 7290 730
rect -312 -1288 -250 -1254
rect -312 -1322 -296 -1288
rect -260 -1322 -250 -1288
rect -312 -1354 -250 -1322
<< nsubdiff >>
rect 7230 1020 7290 1050
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
rect -330 -968 -270 -934
rect -330 -1002 -316 -968
rect -282 -1002 -270 -968
rect -330 -1034 -270 -1002
<< psubdiffcont >>
rect 7240 730 7280 770
rect -296 -1322 -260 -1288
<< nsubdiffcont >>
rect 7240 980 7280 1020
rect -316 -1002 -282 -968
<< locali >>
rect 5980 1540 6080 1560
rect 5980 1500 6010 1540
rect 6050 1500 6080 1540
rect 7230 1020 7290 1050
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7230 700 7290 730
rect -330 -968 -270 -934
rect 240 -960 350 -900
rect -330 -1002 -316 -968
rect -282 -1002 -270 -968
rect -330 -1034 -270 -1002
rect -312 -1288 -250 -1254
rect -312 -1322 -296 -1288
rect -260 -1322 -250 -1288
rect -312 -1354 -250 -1322
<< viali >>
rect 2600 5860 2640 5900
rect 3180 5860 3220 5900
rect 3760 5860 3800 5900
rect 4620 5860 4660 5900
rect 5480 5860 5520 5900
rect 6060 5860 6100 5900
rect 6640 5860 6680 5900
rect 7500 5860 7540 5900
rect 8360 5860 8400 5900
rect 8940 5860 8980 5900
rect 5330 1740 5370 1780
rect 5910 1740 5950 1780
rect 6490 1740 6530 1780
rect 7350 1740 7390 1780
rect 8210 1740 8250 1780
rect 8790 1740 8830 1780
rect 9370 1740 9410 1780
rect 10230 1740 10270 1780
rect 6010 1500 6050 1540
rect 7028 1050 7062 1084
rect 7028 974 7062 1008
rect 7240 980 7280 1020
rect 6846 854 6880 888
rect 7240 730 7280 770
rect -140 -1180 -100 -1140
rect 198 -1178 232 -1144
rect -296 -1322 -260 -1288
<< metal1 >>
rect 7020 1084 7070 1100
rect 7020 1050 7028 1084
rect 7062 1050 7070 1084
rect 7020 1008 7070 1050
rect 7020 974 7028 1008
rect 7062 974 7070 1008
rect 2540 870 2640 960
rect 6760 888 6896 908
rect 2540 770 5590 870
rect 6760 854 6846 888
rect 6880 854 6896 888
rect 7020 900 7070 974
rect 7230 1020 7290 1050
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
rect 7350 900 8270 930
rect 7020 860 8270 900
rect 7037 858 8270 860
rect 6760 836 6896 854
rect 7350 830 8270 858
rect 2540 480 2640 770
rect 3960 480 4060 590
rect 3750 380 4390 480
rect 5490 470 5590 770
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7230 700 7290 730
rect 8170 350 8270 830
rect 11080 -70 11180 -50
rect 11080 -130 11100 -70
rect 11160 -130 11180 -70
rect 11080 -150 11180 -130
rect 11840 -70 11940 -50
rect 11840 -130 11860 -70
rect 11920 -130 11940 -70
rect -330 -1034 -270 -934
rect -180 -1140 -94 -1110
rect -280 -1180 -140 -1140
rect -100 -1180 -94 -1140
rect -280 -1200 -94 -1180
rect 192 -1142 242 -1116
rect 192 -1144 330 -1142
rect 192 -1178 198 -1144
rect 232 -1178 330 -1144
rect 192 -1210 242 -1178
rect -312 -1288 -250 -1254
rect -312 -1322 -296 -1288
rect -260 -1322 -250 -1288
rect -312 -1354 -250 -1322
rect 11840 -1430 11940 -130
rect 8140 -1530 11940 -1430
rect 8140 -1960 8240 -1530
rect 11080 -2410 11180 -2390
rect 11080 -2470 11100 -2410
rect 11160 -2470 11180 -2410
rect 11080 -2500 11180 -2470
<< via1 >>
rect 11100 -130 11160 -70
rect 11860 -130 11920 -70
rect 11100 -2470 11160 -2410
<< metal2 >>
rect 11080 -70 11940 -50
rect 11080 -130 11100 -70
rect 11160 -130 11860 -70
rect 11920 -130 11940 -70
rect 11080 -150 11940 -130
rect 11080 -2410 11890 -2390
rect 11080 -2470 11100 -2410
rect 11160 -2470 11890 -2410
rect 11080 -2490 11890 -2470
use dco_freq  dco_freq_0
timestamp 1726743291
transform 1 0 8320 0 1 50
box -880 -1250 3330 640
use dco_freq  dco_freq_1
timestamp 1726743291
transform 1 0 8320 0 1 -2290
box -880 -1250 3330 640
use dco_idac  dco_idac_0
timestamp 1726728476
transform 1 0 2860 0 1 -60
box -1860 -3160 3220 740
use dco_ring_osc  dco_ring_osc_0
timestamp 1726107115
transform 1 0 1680 0 1 4000
box -500 -2520 9440 2160
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 6808 0 1 638
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -202 0 1 -1392
box -38 -48 498 592
<< labels >>
rlabel locali 6040 1560 6040 1560 1 Isup
rlabel metal1 4010 590 4010 590 1 Vbs_34
rlabel metal1 2590 960 2590 960 1 Vbs_12
rlabel metal2 11900 -50 11900 -50 1 ro_div2
rlabel metal2 11820 -2390 11820 -2390 1 pha_DCO
<< end >>
