** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/ALib_VCO_tb.sch
**.subckt ALib_VCO_tb
VDD VDDA GND DC=1.8
Venb1 ENB GND DC=0 PULSE( 0 1.8 0 0.1n 0.1n 20n 1)
V_input Anlg_in GND DC=0 sin(0.8 0.4 0.5Meg 0 0 0)
x1 VDDA ENB GND GND VDD VDD einvp sky130_fd_sc_hd__einvp_1
Xro_1 V_ctrl VDDA pha_0 pha_1 pha_2 pha_3 pha_4 net1 net2 net3 net4 einvp GND 5s_cc_osc
R3 V_ctrl Anlg_in sky130_fd_pr__res_generic_po W=0.482 L=2 m=1
R1 GND V_ctrl sky130_fd_pr__res_generic_po W=0.482 L=2 m=1
**** begin user architecture code


**LIB with Local Computer
*.lib /home/toind/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
*.inc /home/toind/eda/uniccass/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.lib /home/dkits/openpdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /home/dkits/openpdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice




.control
*save all
set nobreak
set num_threads=10
set mode=1
if ($mode = 1)
    save all
    TRAN 1n 100u
    plot Anlg_in V_ctrl pha_0
    MEAS TRAN prd TRIG pha_0 VAL=0.8 RISE=2 TARG pha_0 VAL=0.8 RISE=8
    let freq=6/prd
    echo "Frequency: "
    print freq
end

if ($mode = 2)
    save "VDD" @Vsup[i] "p[0]"
    TRAN 1n 10u
    MEAS TRAN I_vco AVG @Vsup[i] FROM=2u TO=8u
    MEAS TRAN V_vco AVG VDD FROM=2u TO=8u
    let Power=I_vco*V_vco
    echo "Power: "
    print Power
end
.endc


**** end user architecture code
**.ends

* expanding   symbol:  5s_cc_osc.sym # of pins=13
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/5s_cc_osc.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/5s_cc_osc.sch
.subckt 5s_cc_osc VGND VDDA p[0] p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4] GND
*.iopin VDDA
*.iopin VGND
*.opin pn[0]
*.iopin p[0]
*.opin pn[1]
*.opin p[1]
*.opin p[2]
*.opin p[3]
*.opin p[4]
*.opin pn[2]
*.opin pn[3]
*.opin pn[4]
*.iopin GND
Xi_1 p[4] pn[4] VDDA VGND p[0] pn[0] GND cc_inv
Xi_2 p[0] pn[0] VDDA VGND p[1] pn[1] GND cc_inv
Xi_3 p[1] pn[1] VDDA VGND p[2] pn[2] GND cc_inv
Xi_4 p[2] pn[2] VDDA VGND p[3] pn[3] GND cc_inv
Xi_6 p[3] pn[3] VDDA VGND p[4] pn[4] GND cc_inv
.ends


* expanding   symbol:  cc_inv.sym # of pins=7
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/cc_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/cc_inv.sch
.subckt cc_inv inp inn VDDA VGND outp outn GND
*.opin outp
*.ipin inn
*.iopin VGND
*.opin outn
*.ipin inp
*.iopin VDDA
*.iopin GND
Xi_1 VDDA VGND outp GND inp main_inv
Xi_2 VDDA VGND outn GND inn main_inv
Xi_3 VDDA VGND outn GND outp aux_inv
Xi_4 VDDA VGND outp GND outn aux_inv
.ends


* expanding   symbol:  main_inv.sym # of pins=5
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sch
.subckt main_inv VDDA VGND Y GND A
*.iopin VDDA
*.iopin VGND
*.ipin A
*.opin Y
*.iopin GND
XM1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  aux_inv.sym # of pins=5
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sch
.subckt aux_inv VDDA VGND Y GND A
*.iopin VDDA
*.iopin VGND
*.ipin A
*.opin Y
*.iopin GND
XM1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDDA
.end
