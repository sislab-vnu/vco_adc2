magic
tech sky130A
magscale 1 2
timestamp 1726742472
<< nwell >>
rect -100 0 0 440
rect 1400 0 1500 440
<< poly >>
rect -320 500 -220 520
rect -320 460 -300 500
rect -240 460 -220 500
rect -320 440 -220 460
rect 120 500 580 520
rect 120 460 140 500
rect 180 460 220 500
rect 260 460 300 500
rect 340 460 380 500
rect 420 460 460 500
rect 500 460 580 500
rect 120 440 580 460
rect 820 500 1280 520
rect 820 460 840 500
rect 880 460 920 500
rect 960 460 1000 500
rect 1040 460 1080 500
rect 1120 460 1160 500
rect 1200 460 1280 500
rect 820 440 1280 460
rect 1620 500 1720 520
rect 1620 460 1640 500
rect 1700 460 1720 500
rect 1620 440 1720 460
rect 200 -420 480 -400
rect 200 -460 220 -420
rect 260 -460 320 -420
rect 360 -460 420 -420
rect 460 -460 480 -420
rect 200 -480 480 -460
rect 920 -980 1200 -960
rect 920 -1020 940 -980
rect 980 -1020 1040 -980
rect 1080 -1020 1140 -980
rect 1180 -1020 1200 -980
rect 920 -1040 1200 -1020
rect -640 -1160 -360 -1140
rect -640 -1200 -620 -1160
rect -580 -1200 -520 -1160
rect -480 -1200 -420 -1160
rect -380 -1200 -360 -1160
rect -640 -1220 -360 -1200
rect 1760 -1160 2040 -1140
rect 1760 -1200 1780 -1160
rect 1820 -1200 1880 -1160
rect 1920 -1200 1980 -1160
rect 2020 -1200 2040 -1160
rect 1760 -1220 2040 -1200
rect 610 -1838 690 -1770
<< polycont >>
rect -300 460 -240 500
rect 140 460 180 500
rect 220 460 260 500
rect 300 460 340 500
rect 380 460 420 500
rect 460 460 500 500
rect 840 460 880 500
rect 920 460 960 500
rect 1000 460 1040 500
rect 1080 460 1120 500
rect 1160 460 1200 500
rect 1640 460 1700 500
rect 220 -460 260 -420
rect 320 -460 360 -420
rect 420 -460 460 -420
rect 940 -1020 980 -980
rect 1040 -1020 1080 -980
rect 1140 -1020 1180 -980
rect -620 -1200 -580 -1160
rect -520 -1200 -480 -1160
rect -420 -1200 -380 -1160
rect 1780 -1200 1820 -1160
rect 1880 -1200 1920 -1160
rect 1980 -1200 2020 -1160
<< locali >>
rect -480 660 1540 740
rect -480 320 -400 660
rect -320 500 -220 520
rect -320 460 -300 500
rect -240 460 -220 500
rect -320 440 -220 460
rect 120 500 580 520
rect 120 460 140 500
rect 180 460 220 500
rect 260 460 300 500
rect 340 460 380 500
rect 420 460 460 500
rect 500 460 580 500
rect 120 440 580 460
rect 820 500 1280 520
rect 820 460 840 500
rect 880 460 920 500
rect 960 460 1000 500
rect 1040 460 1080 500
rect 1120 460 1160 500
rect 1200 460 1280 500
rect 820 440 1280 460
rect 1460 340 1540 660
rect 1620 500 1720 520
rect 1620 460 1640 500
rect 1700 460 1720 500
rect 1620 440 1720 460
rect -140 160 40 320
rect 660 160 740 320
rect 1800 40 2120 120
rect 1280 -100 1360 40
rect -720 -180 1760 -100
rect -720 -300 -640 -180
rect 40 -600 120 -180
rect 200 -420 480 -400
rect 200 -460 220 -420
rect 260 -460 320 -420
rect 360 -460 420 -420
rect 460 -460 480 -420
rect 200 -480 480 -460
rect 1280 -600 1360 -180
rect 1680 -300 1760 -180
rect 2040 -300 2120 40
rect 740 -920 840 -840
rect 480 -1030 560 -920
rect -280 -1100 560 -1030
rect -640 -1160 -360 -1140
rect -640 -1200 -620 -1160
rect -580 -1200 -520 -1160
rect -480 -1200 -420 -1160
rect -380 -1200 -360 -1160
rect -640 -1220 -360 -1200
rect -280 -2270 -200 -1100
rect 740 -1300 820 -920
rect 920 -980 1200 -960
rect 920 -1020 940 -980
rect 980 -1020 1040 -980
rect 1080 -1020 1140 -980
rect 1180 -1020 1200 -980
rect 920 -1040 1200 -1020
rect 1760 -1160 2040 -1140
rect 1760 -1200 1780 -1160
rect 1820 -1200 1880 -1160
rect 1920 -1200 1980 -1160
rect 2020 -1200 2040 -1160
rect 1760 -1220 2040 -1200
rect 2120 -1300 2200 -1020
rect 740 -1322 2200 -1300
rect 740 -1356 2146 -1322
rect 2180 -1356 2200 -1322
rect 740 -1380 2200 -1356
rect 610 -1790 690 -1770
rect 440 -1792 1080 -1790
rect 440 -1826 632 -1792
rect 666 -1826 1080 -1792
rect 440 -1830 1080 -1826
rect 1228 -1796 1520 -1792
rect 1228 -1830 1462 -1796
rect 1496 -1830 1520 -1796
rect 610 -1838 690 -1830
rect 1228 -1836 1520 -1830
<< viali >>
rect -300 460 -240 500
rect 140 460 180 500
rect 220 460 260 500
rect 300 460 340 500
rect 380 460 420 500
rect 460 460 500 500
rect 840 460 880 500
rect 920 460 960 500
rect 1000 460 1040 500
rect 1080 460 1120 500
rect 1160 460 1200 500
rect 1640 460 1700 500
rect 220 -460 260 -420
rect 320 -460 360 -420
rect 420 -460 460 -420
rect -620 -1200 -580 -1160
rect -520 -1200 -480 -1160
rect -420 -1200 -380 -1160
rect 940 -1020 980 -980
rect 1040 -1020 1080 -980
rect 1140 -1020 1180 -980
rect 1780 -1200 1820 -1160
rect 1880 -1200 1920 -1160
rect 1980 -1200 2020 -1160
rect 2146 -1356 2180 -1322
rect 216 -1836 250 -1802
rect 632 -1826 666 -1792
rect 1462 -1830 1496 -1796
<< metal1 >>
rect -320 500 -220 840
rect 300 520 400 840
rect 1000 520 1120 840
rect -320 460 -300 500
rect -240 460 -220 500
rect -320 440 -220 460
rect 120 500 580 520
rect 120 460 140 500
rect 180 460 220 500
rect 260 460 300 500
rect 340 460 380 500
rect 420 460 460 500
rect 500 460 580 500
rect 120 440 580 460
rect 820 500 1280 520
rect 820 460 840 500
rect 880 460 920 500
rect 960 460 1000 500
rect 1040 460 1080 500
rect 1120 460 1160 500
rect 1200 460 1280 500
rect 820 440 1280 460
rect 1620 500 1720 840
rect 1620 460 1640 500
rect 1700 460 1720 500
rect 1620 440 1720 460
rect 300 -360 1520 -280
rect 300 -400 380 -360
rect 200 -420 480 -400
rect 200 -460 220 -420
rect 260 -460 320 -420
rect 360 -460 420 -420
rect 460 -460 480 -420
rect 200 -480 480 -460
rect 610 -980 1200 -960
rect 610 -1020 940 -980
rect 980 -1020 1040 -980
rect 1080 -1020 1140 -980
rect 1180 -1020 1200 -980
rect 610 -1040 1200 -1020
rect 610 -1140 690 -1040
rect -640 -1160 690 -1140
rect -640 -1200 -620 -1160
rect -580 -1200 -520 -1160
rect -480 -1200 -420 -1160
rect -380 -1200 690 -1160
rect -640 -1220 690 -1200
rect 2 -1802 266 -1782
rect 2 -1836 216 -1802
rect 250 -1836 266 -1802
rect 2 -1854 266 -1836
rect 610 -1792 690 -1220
rect 610 -1826 632 -1792
rect 666 -1826 690 -1792
rect 610 -1838 690 -1826
rect 1440 -1140 1520 -360
rect 1440 -1160 2040 -1140
rect 1440 -1200 1780 -1160
rect 1820 -1200 1880 -1160
rect 1920 -1200 1980 -1160
rect 2020 -1200 2040 -1160
rect 1440 -1220 2040 -1200
rect 1440 -1796 1520 -1220
rect 2120 -1322 2326 -1300
rect 2120 -1356 2146 -1322
rect 2180 -1356 2326 -1322
rect 2120 -1380 2326 -1356
rect 1440 -1830 1462 -1796
rect 1496 -1830 1520 -1796
rect 1440 -1836 1520 -1830
use nmos_idac_lk  nmos_idac_lk_0
timestamp 1723695905
transform 1 0 200 0 1 -920
box -120 -40 400 440
use nmos_idac_lk  nmos_idac_lk_1
timestamp 1723695905
transform 1 0 920 0 1 -920
box -120 -40 400 440
use pmos_idac_br2  pmos_idac_br2_0
timestamp 1723704601
transform 1 0 120 0 1 40
box -120 -40 580 400
use pmos_idac_br2  pmos_idac_br2_1
timestamp 1723704601
transform 1 0 820 0 1 40
box -120 -40 580 400
use pmos_idac_br  pmos_idac_br_0
timestamp 1723711581
transform 1 0 -320 0 1 40
box -120 -40 220 400
use pmos_idac_br  pmos_idac_br_1
timestamp 1723711581
transform 1 0 1620 0 1 40
box -120 -40 220 400
use pmos_idac_lk  pmos_idac_lk_0
timestamp 1723695758
transform 1 0 -640 0 1 -1100
box -120 -40 400 840
use pmos_idac_lk  pmos_idac_lk_1
timestamp 1723695758
transform 1 0 1760 0 1 -1100
box -120 -40 400 840
use sky130_fd_pr__res_xhigh_po_0p35_JPCEFB  sky130_fd_pr__res_xhigh_po_0p35_JPCEFB_0
timestamp 1723776395
transform 0 1 772 -1 0 -2305
box -35 -1272 35 1272
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 178 0 1 -2052
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 1058 0 1 -2052
box -38 -48 314 592
<< end >>
