* NGSPICE file created from vco_adc2.ext - technology: sky130A

.subckt aux_inv A Y VGND VDDA GND
X0 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt main_inv A Y VGND GND VDDA
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt cc_inv inp inn outp outn VGND GND VDDA
Xaux_inv_0 outp outn VGND VDDA GND aux_inv
Xaux_inv_1 outn outp VGND VDDA GND aux_inv
Xmain_inv_0 inp outp VGND GND VDDA main_inv
Xmain_inv_1 inn outn VGND GND VDDA main_inv
.ends

.subckt x5s_cc_osc pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VGND VDDA
+ GND
Xcc_inv_0 p[4] pn[4] p[0] pn[0] VGND GND VDDA cc_inv
Xcc_inv_1 p[0] pn[0] p[1] pn[1] VGND GND VDDA cc_inv
Xcc_inv_2 p[1] pn[1] p[2] pn[2] VGND GND VDDA cc_inv
Xcc_inv_3 p[3] pn[3] p[4] pn[4] VGND GND VDDA cc_inv
Xcc_inv_4 p[2] pn[2] p[3] pn[3] VGND GND VDDA cc_inv
.ends

.subckt sky130_fd_pr__res_generic_po_DKCPUZ a_n48_200# a_n48_n630#
R0 a_n48_200# a_n48_n630# sky130_fd_pr__res_generic_po w=0.48 l=2
.ends


.subckt ALib_VCO Anlg_in ENB GND p[4] VDDA
Xx5s_cc_osc_0 x5s_cc_osc_0/pn[0] x5s_cc_osc_0/pn[1] x5s_cc_osc_0/pn[2] x5s_cc_osc_0/pn[3]
+ pn[4] x5s_cc_osc_0/p[0] x5s_cc_osc_0/p[1] x5s_cc_osc_0/p[2] x5s_cc_osc_0/p[3] p[4]
+ Vctrl VDDA GND x5s_cc_osc
Xsky130_fd_pr__res_generic_po_DKCPUZ_0 Vctrl Anlg_in sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_pr__res_generic_po_DKCPUZ_1 Vctrl GND sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_sc_hd__einvp_1_0 VDDA ENB GND GND VDDA VDDA pn[4] sky130_fd_sc_hd__einvp_1
.ends






.subckt DLib_Quantizer D CLK Dout FBack VDDA GND
Xsky130_fd_sc_hd__dlygate4sd3_1_0 CLK GND GND VDDA VDDA DL1 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_1 DL1 GND GND VDDA VDDA DL2 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__inv_2_0 FBack_inv GND GND VDDA VDDA FBack sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_0 D GND GND VDDA VDDA sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dlygate4sd3_1_2 DL2 GND GND VDDA VDDA DL3 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_3 DL3 GND GND VDDA VDDA DL4 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_4 DL4 GND GND VDDA VDDA DL5 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_5 DL5 GND GND VDDA VDDA CLK_dly sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__nand2_1_0 CLK_dly Dout GND GND VDDA VDDA FBack_inv sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_0 CLK sky130_fd_sc_hd__buf_2_0/X GND GND VDDA VDDA Dout
+ sky130_fd_sc_hd__dfxtp_1
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_RSCMUS a_n35_n1272# a_n35_840# a_n165_n1402#
X0 a_n35_840# a_n35_n1272# a_n165_n1402# sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

.subckt ALib_IDAC Vbs1 Vbs2 Vbs3 Vbs4 Dctrl Isup VDDA GND
Xsky130_fd_sc_hd__buf_2_0 Dctrl GND GND VDDA VDDA sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A GND GND VDDA VDDA sky130_fd_sc_hd__inv_2_0/Y
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0 GND a_n150_n1850# GND sky130_fd_pr__res_xhigh_po_0p35_RSCMUS
X0 Isup sky130_fd_sc_hd__inv_2_0/A w_n510_n1930# GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X1 w_2370_n90# Vbs1 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X2 w_n510_n1930# Vbs4 w_1270_n80# w_1270_n80# sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X3 a_n150_n1850# sky130_fd_sc_hd__inv_2_0/Y w_n510_n1930# GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X4 Isup sky130_fd_sc_hd__inv_2_0/Y w_n510_n1930# w_n510_n1930# sky130_fd_pr__pfet_01v8_hvt ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
X5 w_1270_n80# Vbs3 VDDA VDDA sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X6 Isup Vbs2 w_2370_n90# w_2370_n90# sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X7 w_n510_n1930# sky130_fd_sc_hd__inv_2_0/A a_n150_n1850# w_n510_n1930# sky130_fd_pr__pfet_01v8_hvt ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.5 M=2
.ends




.subckt DLib_freqDiv2 clk clkDiv2 VDDA GND
Xsky130_fd_sc_hd__buf_4_0 Q_N GND GND VDDA VDDA Q_N_buf sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_4_0 clk GND GND VDDA VDDA clkinv sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__dfxtp_1_0 clkinv Q_N_buf GND GND VDDA VDDA D sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxbp_2_0 clk D GND GND VDDA VDDA clkDiv2 Q_N sky130_fd_sc_hd__dfxbp_2
.ends

.subckt aux_inv_dco A Y VDDA VGND
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.2
X1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=1.2
.ends

.subckt main_inv_dco A Y VDDA VGND
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=1.2 M=2
X1 VGND A Y VGND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=1.2 M=2
.ends

.subckt cc_inv_dco outp outn VDDA inn inp VGND
Xaux_inv_dco_0 outp outn VDDA VGND aux_inv_dco
Xaux_inv_dco_1 outn outp VDDA VGND aux_inv_dco
Xmain_inv_dco_0 inp outp VDDA VGND main_inv_dco
Xmain_inv_dco_1 inn outn VDDA VGND main_inv_dco
.ends

.subckt x5s_cc_osc_dco pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VDDA
+ VGND
Xcc_inv_dco_1 p[1] pn[1] VDDA pn[0] p[0] VGND cc_inv_dco
Xcc_inv_dco_2 p[2] pn[2] VDDA pn[1] p[1] VGND cc_inv_dco
Xcc_inv_dco_3 p[4] pn[4] VDDA pn[3] p[3] VGND cc_inv_dco
Xcc_inv_dco_4 p[3] pn[3] VDDA pn[2] p[2] VGND cc_inv_dco
Xcc_inv_dco_0 p[0] pn[0] VDDA pn[4] p[4] VGND cc_inv_dco
.ends

.subckt ALib_DCO Vbs_12 Vbs_34 pha_DCO Dctrl ENB VDDA GND
Xsky130_fd_sc_hd__buf_2_0 x5s_cc_osc_dco_0/p[4] GND GND VDDA VDDA DLib_freqDiv2_1/clk
+ sky130_fd_sc_hd__buf_2
XALib_IDAC_0 Vbs_12 Vbs_12 Vbs_34 Vbs_34 Dctrl ALib_IDAC_0/Isup VDDA GND ALib_IDAC
XDLib_freqDiv2_0 DLib_freqDiv2_0/clk pha_DCO VDDA GND DLib_freqDiv2
XDLib_freqDiv2_1 DLib_freqDiv2_1/clk DLib_freqDiv2_0/clk VDDA GND DLib_freqDiv2
Xx5s_cc_osc_dco_0 x5s_cc_osc_dco_0/pn[0] x5s_cc_osc_dco_0/pn[1] x5s_cc_osc_dco_0/pn[2]
+ x5s_cc_osc_dco_0/pn[3] x5s_cc_osc_dco_0/pn[4] x5s_cc_osc_dco_0/p[0] x5s_cc_osc_dco_0/p[1]
+ x5s_cc_osc_dco_0/p[2] x5s_cc_osc_dco_0/p[3] x5s_cc_osc_dco_0/p[4] ALib_IDAC_0/Isup
+ GND x5s_cc_osc_dco
Xsky130_fd_sc_hd__einvp_1_0 VDDA ENB GND GND VDDA VDDA x5s_cc_osc_dco_0/pn[4] sky130_fd_sc_hd__einvp_1
.ends



.subckt DLib_UpDownCounter UP DOWN setB VDDA GND Dout_buf
Xsky130_fd_sc_hd__dfstp_1_0 UP_buf Q2N SetBi GND GND VDDA VDDA Q1 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfstp_1_1 DWN_buf Q1_buf SetBi GND GND VDDA VDDA Q2 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__inv_2_0 setB GND GND VDDA VDDA SetBi sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_1 DOWN GND GND VDDA VDDA DWN_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_1 Q2 GND GND VDDA VDDA Q2N sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_2 Dout GND GND VDDA VDDA Dout_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_3 Q1 GND GND VDDA VDDA Q1_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_4 UP GND GND VDDA VDDA UP_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_1 Q1 Q2 GND GND VDDA VDDA Dout sky130_fd_sc_hd__xor2_1
.ends

.subckt vco_adc2 vbias_12 vbias_34 analog_in enable_in clk quantizer_out VDDA GND
XALib_VCO_0 analog_in enable_in GND ALib_VCO_0/p[4] VDDA ALib_VCO
XDLib_Quantizer_0 DLib_Quantizer_0/D clk quantizer_out DLib_Quantizer_0/FBack VDDA
+ GND DLib_Quantizer
XALib_DCO_0 vbias_12 vbias_34 ALib_DCO_0/pha_DCO ALib_DCO_0/Dctrl enable_in VDDA GND
+ ALib_DCO
XDLib_UpDownCounter_0 ALib_DCO_0/pha_DCO DLib_Quantizer_0/FBack enable_in VDDA GND
+ DLib_Quantizer_0/D DLib_UpDownCounter
XDLib_UpDownCounter_1 ALib_VCO_0/p[4] DLib_Quantizer_0/FBack enable_in VDDA GND ALib_DCO_0/Dctrl
+ DLib_UpDownCounter
.ends


