magic
tech sky130A
magscale 1 2
timestamp 1727087206
<< nwell >>
rect -860 -780 2690 -440
rect -850 -1500 -670 -1480
rect -850 -1810 -690 -1500
rect -850 -1820 -680 -1810
rect 1610 -1910 1810 -1580
rect -190 -2840 -20 -2820
rect 1960 -2830 2320 -2820
rect -190 -3140 -40 -2840
rect 1960 -3140 2280 -2830
rect -190 -3150 -20 -3140
rect 1960 -3150 2350 -3140
<< pwell >>
rect -860 -1010 -690 -870
rect -390 -1010 -10 -870
rect 1840 -1010 2290 -870
rect -850 -2050 -660 -1870
rect 1570 -2150 1850 -2010
rect -230 -2770 70 -2580
rect 1920 -2720 2320 -2580
<< psubdiff >>
rect -820 -910 -740 -880
rect -820 -950 -800 -910
rect -760 -950 -740 -910
rect -820 -980 -740 -950
rect -810 -1950 -730 -1920
rect -810 -1990 -790 -1950
rect -750 -1990 -730 -1950
rect -810 -2020 -730 -1990
rect 1660 -2060 1760 -2040
rect 1660 -2100 1690 -2060
rect 1730 -2100 1760 -2060
rect 1660 -2120 1760 -2100
rect 2140 -2630 2240 -2610
rect 2140 -2670 2170 -2630
rect 2210 -2670 2240 -2630
rect 2140 -2690 2240 -2670
<< nsubdiff >>
rect -210 -590 -130 -560
rect -210 -630 -190 -590
rect -150 -630 -130 -590
rect -210 -660 -130 -630
rect -810 -1600 -730 -1570
rect -810 -1640 -790 -1600
rect -750 -1640 -730 -1600
rect -810 -1670 -730 -1640
rect 1680 -1750 1760 -1720
rect 1680 -1790 1700 -1750
rect 1740 -1790 1760 -1750
rect 1680 -1820 1760 -1790
rect -130 -2940 -50 -2910
rect -130 -2980 -110 -2940
rect -70 -2980 -50 -2940
rect -130 -3010 -50 -2980
<< psubdiffcont >>
rect -800 -950 -760 -910
rect -790 -1990 -750 -1950
rect 1690 -2100 1730 -2060
rect 2170 -2670 2210 -2630
<< nsubdiffcont >>
rect -190 -630 -150 -590
rect -790 -1640 -750 -1600
rect 1700 -1790 1740 -1750
rect -110 -2980 -70 -2940
<< locali >>
rect 2630 -540 3140 -470
rect -210 -590 -130 -560
rect -210 -630 -190 -590
rect -150 -630 -130 -590
rect -210 -660 -130 -630
rect -880 -830 -610 -760
rect -440 -810 20 -770
rect 1820 -780 2300 -760
rect 1820 -820 2100 -780
rect 2140 -820 2300 -780
rect 1820 -840 2300 -820
rect -820 -910 -740 -880
rect -820 -950 -800 -910
rect -760 -950 -740 -910
rect -820 -980 -740 -950
rect -360 -1080 -10 -980
rect 1910 -1080 2280 -990
rect -810 -1600 -730 -1570
rect -430 -1580 1000 -1510
rect -810 -1640 -790 -1600
rect -750 -1640 -730 -1600
rect 930 -1620 1000 -1580
rect 3070 -1610 3140 -540
rect -810 -1670 -730 -1640
rect 2190 -1680 3140 -1610
rect 1680 -1750 1760 -1720
rect 1680 -1790 1700 -1750
rect 1740 -1790 1760 -1750
rect 1680 -1820 1760 -1790
rect 1460 -1900 1800 -1890
rect -810 -1950 -730 -1920
rect -810 -1990 -790 -1950
rect -750 -1990 -730 -1950
rect 1460 -1940 1870 -1900
rect 2090 -1950 2100 -1940
rect -810 -2020 -730 -1990
rect -430 -2030 510 -2020
rect -430 -2070 450 -2030
rect 490 -2070 510 -2030
rect -430 -2090 510 -2070
rect 440 -2130 510 -2090
rect 1660 -2060 1760 -2040
rect 1660 -2100 1690 -2060
rect 1730 -2100 1760 -2060
rect 1660 -2120 1760 -2100
rect 440 -2200 970 -2130
rect -250 -2610 10 -2520
rect 440 -2565 510 -2200
rect 1920 -2610 2350 -2540
rect 2140 -2630 2240 -2610
rect 2140 -2670 2170 -2630
rect 2210 -2670 2240 -2630
rect 2140 -2690 2240 -2670
rect 2720 -2758 2830 -2750
rect 1870 -2770 2220 -2760
rect -248 -2826 106 -2778
rect 1870 -2810 2170 -2770
rect 2210 -2810 2220 -2770
rect 1880 -2830 2220 -2810
rect 2592 -2834 2830 -2758
rect 2720 -2840 2830 -2834
rect -130 -2940 -50 -2910
rect -130 -2980 -110 -2940
rect -70 -2980 -50 -2940
rect -130 -3010 -50 -2980
rect 3070 -3080 3140 -1680
rect 2670 -3150 3140 -3080
<< viali >>
rect -190 -630 -150 -590
rect 2502 -662 2536 -628
rect 360 -790 400 -750
rect 2100 -820 2140 -780
rect -800 -950 -760 -910
rect -790 -1640 -750 -1600
rect 1700 -1790 1740 -1750
rect -638 -1854 -598 -1814
rect 2064 -1810 2104 -1770
rect -534 -1854 -500 -1820
rect -790 -1990 -750 -1950
rect 1024 -1952 1058 -1918
rect 1138 -1950 1172 -1916
rect 450 -2070 490 -2030
rect 1690 -2100 1730 -2060
rect 2170 -2670 2210 -2630
rect -386 -2726 -346 -2686
rect 92 -2714 132 -2674
rect 2170 -2810 2210 -2770
rect 1520 -2850 1560 -2810
rect -110 -2980 -70 -2940
rect 2424 -2942 2458 -2908
<< metal1 >>
rect -690 -530 -680 -440
rect -340 -540 0 -440
rect 1910 -540 2280 -440
rect -210 -590 -130 -540
rect -210 -630 -190 -590
rect -150 -630 -130 -590
rect -210 -660 -130 -630
rect 2490 -628 2950 -610
rect 2490 -662 2502 -628
rect 2536 -662 2950 -628
rect 2490 -680 2950 -662
rect -210 -750 420 -730
rect -210 -790 360 -750
rect 400 -790 420 -750
rect -210 -810 420 -790
rect 2080 -780 2150 -760
rect -820 -910 -740 -880
rect -820 -950 -800 -910
rect -760 -950 -740 -910
rect -820 -980 -740 -950
rect -820 -1080 -680 -980
rect -810 -1580 -660 -1480
rect -810 -1600 -730 -1580
rect -810 -1640 -790 -1600
rect -750 -1640 -730 -1600
rect -810 -1670 -730 -1640
rect -470 -1800 -380 -1790
rect -830 -1814 -580 -1800
rect -830 -1854 -638 -1814
rect -598 -1854 -580 -1814
rect -830 -1870 -580 -1854
rect -550 -1820 -450 -1800
rect -550 -1854 -534 -1820
rect -500 -1854 -450 -1820
rect -550 -1860 -450 -1854
rect -390 -1860 -380 -1800
rect -550 -1870 -380 -1860
rect -470 -1880 -380 -1870
rect -810 -1950 -730 -1920
rect -810 -1990 -790 -1950
rect -750 -1990 -730 -1950
rect -810 -2020 -730 -1990
rect -810 -2130 -670 -2020
rect -210 -2180 -140 -810
rect 2080 -820 2100 -780
rect 2140 -820 2150 -780
rect 730 -860 830 -840
rect 730 -920 750 -860
rect 810 -920 830 -860
rect 730 -930 830 -920
rect 440 -2030 510 -1070
rect 2080 -1330 2150 -820
rect 610 -1400 2150 -1330
rect 610 -1730 680 -1400
rect 1570 -1670 1850 -1570
rect 610 -1800 1190 -1730
rect 1000 -1918 1070 -1900
rect 1120 -1910 1190 -1800
rect 1680 -1750 1760 -1670
rect 1680 -1790 1700 -1750
rect 1740 -1790 1760 -1750
rect 1680 -1820 1760 -1790
rect 2050 -1770 2110 -1750
rect 2050 -1810 2064 -1770
rect 2104 -1810 2110 -1770
rect 2050 -1890 2110 -1810
rect 1000 -1952 1024 -1918
rect 1058 -1952 1070 -1918
rect 1000 -1970 1070 -1952
rect 1100 -1916 1210 -1910
rect 1100 -1950 1138 -1916
rect 1172 -1950 1210 -1916
rect 1100 -1960 1210 -1950
rect 2050 -1960 2280 -1890
rect 2050 -1962 2110 -1960
rect 440 -2070 450 -2030
rect 490 -2070 510 -2030
rect 440 -2090 510 -2070
rect 610 -2040 1070 -1970
rect -740 -2240 -140 -2180
rect -740 -2670 -670 -2240
rect 610 -2380 680 -2040
rect 1660 -2060 1760 -2040
rect 1660 -2100 1690 -2060
rect 1730 -2100 1760 -2060
rect 1660 -2120 1760 -2100
rect 1570 -2220 1850 -2120
rect 2880 -2340 2950 -680
rect -140 -2450 680 -2380
rect 2010 -2410 2950 -2340
rect -140 -2660 -70 -2450
rect -740 -2686 -330 -2670
rect -740 -2726 -386 -2686
rect -346 -2726 -330 -2686
rect -740 -2740 -330 -2726
rect -140 -2674 150 -2660
rect -140 -2714 92 -2674
rect 132 -2714 150 -2674
rect -140 -2740 150 -2714
rect 1110 -2670 1210 -2650
rect 1110 -2730 1130 -2670
rect 1190 -2730 1210 -2670
rect 1110 -2750 1210 -2730
rect 1490 -2810 1570 -2780
rect 1490 -2850 1520 -2810
rect 1560 -2820 1570 -2810
rect 2010 -2820 2080 -2410
rect 2140 -2630 2240 -2610
rect 2140 -2670 2170 -2630
rect 2210 -2670 2240 -2630
rect 2140 -2690 2240 -2670
rect 1560 -2850 2080 -2820
rect 2150 -2770 2480 -2760
rect 2150 -2810 2170 -2770
rect 2210 -2810 2480 -2770
rect 2150 -2830 2480 -2810
rect 1490 -2880 2080 -2850
rect 1490 -2890 1730 -2880
rect 1850 -2890 2080 -2880
rect 2410 -2908 2480 -2830
rect -130 -2940 -50 -2910
rect -130 -2980 -110 -2940
rect -70 -2980 -50 -2940
rect -130 -3060 -50 -2980
rect 2410 -2942 2424 -2908
rect 2458 -2942 2480 -2908
rect 2410 -2990 2480 -2942
rect -230 -3150 10 -3060
rect 1920 -3150 2320 -3060
<< via1 >>
rect -450 -1860 -390 -1800
rect 750 -920 810 -860
rect 1130 -2730 1190 -2670
<< metal2 >>
rect 730 -860 830 -840
rect 730 -920 750 -860
rect 810 -920 830 -860
rect 730 -950 830 -920
rect 730 -1180 800 -950
rect 100 -1250 800 -1180
rect -470 -1800 -380 -1790
rect 100 -1800 170 -1250
rect -470 -1860 -450 -1800
rect -390 -1860 170 -1800
rect -470 -1870 170 -1860
rect -470 -1880 -380 -1870
rect 100 -2260 170 -1870
rect 100 -2330 1180 -2260
rect 1110 -2650 1180 -2330
rect 1110 -2670 1210 -2650
rect 1110 -2730 1130 -2670
rect 1190 -2730 1210 -2670
rect 1110 -2750 1210 -2730
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform -1 0 2680 0 -1 -2562
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1709947739
transform 1 0 1846 0 1 -2168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1709947739
transform 1 0 2280 0 1 -1032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_4
timestamp 1709947739
transform 1 0 -702 0 1 -1032
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -14 0 1 -1032
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_1
timestamp 1709947739
transform -1 0 1926 0 -1 -2562
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -672 0 1 -2074
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1709947739
transform -1 0 -224 0 -1 -2562
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 930 0 1 -2168
box -38 -48 682 592
<< labels >>
rlabel locali 2780 -2750 2780 -2750 1 DOWN
port 3 n
rlabel metal1 2770 -610 2770 -610 1 Q1_buf
rlabel locali 2040 -840 2040 -840 5 Q1
rlabel locali 1620 -1940 1620 -1940 5 Dout
rlabel metal1 2270 -1890 2270 -1890 1 Dout_buf
port 4 n
rlabel metal1 850 -1970 850 -1970 1 Q2
rlabel metal1 -780 -1800 -780 -1800 1 SetB
port 2 n
rlabel metal1 -210 -1140 -210 -1140 7 Q2N
rlabel metal2 -330 -1800 -330 -1800 1 SetBi
rlabel locali -280 -810 -280 -810 5 UP_buf
rlabel locali -770 -760 -770 -760 1 UP
port 1 n
rlabel locali -330 -2020 -330 -2020 1 GND
rlabel metal1 2260 -2760 2260 -2760 1 DWN_buf
rlabel locali 2790 -470 2790 -470 1 VCCD
<< end >>
