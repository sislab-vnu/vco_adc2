* NGSPICE file created from x5s_cc_osc_dco.ext - technology: sky130A

.subckt aux_inv_dco A Y VDDA VGND
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.2
X1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=1.2
.ends

.subckt main_inv_dco A Y VDDA VGND
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=1.2 M=2
X1 VGND A Y VGND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=1.2 M=2
.ends

.subckt cc_inv_dco outp outn VDDA inn inp VGND
Xaux_inv_dco_0 outp outn VDDA VGND aux_inv_dco
Xaux_inv_dco_1 outn outp VDDA VGND aux_inv_dco
Xmain_inv_dco_0 inp outp VDDA VGND main_inv_dco
Xmain_inv_dco_1 inn outn VDDA VGND main_inv_dco
.ends

.subckt x5s_cc_osc_dco pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VDDA
+ VGND
Xcc_inv_dco_1 p[1] pn[1] VDDA pn[0] p[0] VGND cc_inv_dco
Xcc_inv_dco_2 p[2] pn[2] VDDA pn[1] p[1] VGND cc_inv_dco
Xcc_inv_dco_3 p[4] pn[4] VDDA pn[3] p[3] VGND cc_inv_dco
Xcc_inv_dco_4 p[3] pn[3] VDDA pn[2] p[2] VGND cc_inv_dco
Xcc_inv_dco_0 p[0] pn[0] VDDA pn[4] p[4] VGND cc_inv_dco
.ends


