magic
tech sky130A
magscale 1 2
timestamp 1731468405
<< nwell >>
rect -580 -80 -100 440
rect 170 -80 1010 440
rect 1270 -80 2110 440
rect 2370 -90 2850 430
rect -1560 -2110 -1230 -1880
rect -510 -1930 150 -970
rect 2260 -1940 2920 -980
<< pwell >>
rect -1790 -2160 -1610 -1850
rect 450 -1560 1110 -1000
rect 1360 -1560 2020 -1000
rect 2630 -2830 2670 -2790
rect 2510 -3090 2650 -2920
<< nmos >>
rect 710 -1480 810 -1080
rect 890 -1480 990 -1080
rect 1480 -1480 1580 -1080
rect 1660 -1480 1760 -1080
<< pmoshvt >>
rect -320 0 -220 360
rect 430 0 530 360
rect 610 0 710 360
rect 790 0 890 360
rect 1530 0 1630 360
rect 1710 0 1810 360
rect 1890 0 1990 360
rect 2630 -10 2730 350
rect -250 -1850 -150 -1050
rect -70 -1850 30 -1050
rect 2520 -1860 2620 -1060
rect 2700 -1860 2800 -1060
<< ndiff >>
rect 630 -1110 710 -1080
rect 630 -1150 650 -1110
rect 690 -1150 710 -1110
rect 630 -1190 710 -1150
rect 630 -1230 650 -1190
rect 690 -1230 710 -1190
rect 630 -1270 710 -1230
rect 630 -1310 650 -1270
rect 690 -1310 710 -1270
rect 630 -1350 710 -1310
rect 630 -1390 650 -1350
rect 690 -1390 710 -1350
rect 630 -1480 710 -1390
rect 810 -1110 890 -1080
rect 810 -1150 830 -1110
rect 870 -1150 890 -1110
rect 810 -1190 890 -1150
rect 810 -1230 830 -1190
rect 870 -1230 890 -1190
rect 810 -1270 890 -1230
rect 810 -1310 830 -1270
rect 870 -1310 890 -1270
rect 810 -1350 890 -1310
rect 810 -1390 830 -1350
rect 870 -1390 890 -1350
rect 810 -1480 890 -1390
rect 990 -1110 1070 -1080
rect 990 -1150 1010 -1110
rect 1050 -1150 1070 -1110
rect 990 -1190 1070 -1150
rect 990 -1230 1010 -1190
rect 1050 -1230 1070 -1190
rect 990 -1270 1070 -1230
rect 990 -1310 1010 -1270
rect 1050 -1310 1070 -1270
rect 990 -1350 1070 -1310
rect 990 -1390 1010 -1350
rect 1050 -1390 1070 -1350
rect 990 -1480 1070 -1390
rect 1400 -1170 1480 -1080
rect 1400 -1210 1420 -1170
rect 1460 -1210 1480 -1170
rect 1400 -1250 1480 -1210
rect 1400 -1290 1420 -1250
rect 1460 -1290 1480 -1250
rect 1400 -1330 1480 -1290
rect 1400 -1370 1420 -1330
rect 1460 -1370 1480 -1330
rect 1400 -1410 1480 -1370
rect 1400 -1450 1420 -1410
rect 1460 -1450 1480 -1410
rect 1400 -1480 1480 -1450
rect 1580 -1170 1660 -1080
rect 1580 -1210 1600 -1170
rect 1640 -1210 1660 -1170
rect 1580 -1250 1660 -1210
rect 1580 -1290 1600 -1250
rect 1640 -1290 1660 -1250
rect 1580 -1330 1660 -1290
rect 1580 -1370 1600 -1330
rect 1640 -1370 1660 -1330
rect 1580 -1410 1660 -1370
rect 1580 -1450 1600 -1410
rect 1640 -1450 1660 -1410
rect 1580 -1480 1660 -1450
rect 1760 -1170 1840 -1080
rect 1760 -1210 1780 -1170
rect 1820 -1210 1840 -1170
rect 1760 -1250 1840 -1210
rect 1760 -1290 1780 -1250
rect 1820 -1290 1840 -1250
rect 1760 -1330 1840 -1290
rect 1760 -1370 1780 -1330
rect 1820 -1370 1840 -1330
rect 1760 -1410 1840 -1370
rect 1760 -1450 1780 -1410
rect 1820 -1450 1840 -1410
rect 1760 -1480 1840 -1450
<< pdiff >>
rect -400 340 -320 360
rect -400 300 -380 340
rect -340 300 -320 340
rect -400 260 -320 300
rect -400 220 -380 260
rect -340 220 -320 260
rect -400 180 -320 220
rect -400 140 -380 180
rect -340 140 -320 180
rect -400 100 -320 140
rect -400 60 -380 100
rect -340 60 -320 100
rect -400 0 -320 60
rect -220 340 -140 360
rect -220 300 -200 340
rect -160 300 -140 340
rect -220 260 -140 300
rect 350 340 430 360
rect 350 300 370 340
rect 410 300 430 340
rect -220 220 -200 260
rect -160 220 -140 260
rect -220 180 -140 220
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 0 -140 60
rect 350 260 430 300
rect 350 220 370 260
rect 410 220 430 260
rect 350 180 430 220
rect 350 140 370 180
rect 410 140 430 180
rect 350 100 430 140
rect 350 60 370 100
rect 410 60 430 100
rect 350 0 430 60
rect 530 340 610 360
rect 530 300 550 340
rect 590 300 610 340
rect 530 260 610 300
rect 530 220 550 260
rect 590 220 610 260
rect 530 180 610 220
rect 530 140 550 180
rect 590 140 610 180
rect 530 100 610 140
rect 530 60 550 100
rect 590 60 610 100
rect 530 0 610 60
rect 710 340 790 360
rect 710 300 730 340
rect 770 300 790 340
rect 710 260 790 300
rect 710 220 730 260
rect 770 220 790 260
rect 710 180 790 220
rect 710 140 730 180
rect 770 140 790 180
rect 710 100 790 140
rect 710 60 730 100
rect 770 60 790 100
rect 710 0 790 60
rect 890 340 970 360
rect 890 300 910 340
rect 950 300 970 340
rect 890 260 970 300
rect 1450 340 1530 360
rect 1450 300 1470 340
rect 1510 300 1530 340
rect 890 220 910 260
rect 950 220 970 260
rect 890 180 970 220
rect 890 140 910 180
rect 950 140 970 180
rect 890 100 970 140
rect 890 60 910 100
rect 950 60 970 100
rect 890 0 970 60
rect 1450 260 1530 300
rect 1450 220 1470 260
rect 1510 220 1530 260
rect 1450 180 1530 220
rect 1450 140 1470 180
rect 1510 140 1530 180
rect 1450 100 1530 140
rect 1450 60 1470 100
rect 1510 60 1530 100
rect 1450 0 1530 60
rect 1630 340 1710 360
rect 1630 300 1650 340
rect 1690 300 1710 340
rect 1630 260 1710 300
rect 1630 220 1650 260
rect 1690 220 1710 260
rect 1630 180 1710 220
rect 1630 140 1650 180
rect 1690 140 1710 180
rect 1630 100 1710 140
rect 1630 60 1650 100
rect 1690 60 1710 100
rect 1630 0 1710 60
rect 1810 340 1890 360
rect 1810 300 1830 340
rect 1870 300 1890 340
rect 1810 260 1890 300
rect 1810 220 1830 260
rect 1870 220 1890 260
rect 1810 180 1890 220
rect 1810 140 1830 180
rect 1870 140 1890 180
rect 1810 100 1890 140
rect 1810 60 1830 100
rect 1870 60 1890 100
rect 1810 0 1890 60
rect 1990 340 2070 360
rect 1990 300 2010 340
rect 2050 300 2070 340
rect 1990 260 2070 300
rect 2550 330 2630 350
rect 2550 290 2570 330
rect 2610 290 2630 330
rect 1990 220 2010 260
rect 2050 220 2070 260
rect 1990 180 2070 220
rect 1990 140 2010 180
rect 2050 140 2070 180
rect 1990 100 2070 140
rect 1990 60 2010 100
rect 2050 60 2070 100
rect 1990 0 2070 60
rect 2550 250 2630 290
rect 2550 210 2570 250
rect 2610 210 2630 250
rect 2550 170 2630 210
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -10 2630 50
rect 2730 330 2810 350
rect 2730 290 2750 330
rect 2790 290 2810 330
rect 2730 250 2810 290
rect 2730 210 2750 250
rect 2790 210 2810 250
rect 2730 170 2810 210
rect 2730 130 2750 170
rect 2790 130 2810 170
rect 2730 90 2810 130
rect 2730 50 2750 90
rect 2790 50 2810 90
rect 2730 -10 2810 50
rect -330 -1070 -250 -1050
rect -330 -1110 -310 -1070
rect -270 -1110 -250 -1070
rect -330 -1150 -250 -1110
rect -330 -1190 -310 -1150
rect -270 -1190 -250 -1150
rect -330 -1230 -250 -1190
rect -330 -1270 -310 -1230
rect -270 -1270 -250 -1230
rect -330 -1310 -250 -1270
rect -330 -1350 -310 -1310
rect -270 -1350 -250 -1310
rect -330 -1390 -250 -1350
rect -330 -1430 -310 -1390
rect -270 -1430 -250 -1390
rect -330 -1470 -250 -1430
rect -330 -1510 -310 -1470
rect -270 -1510 -250 -1470
rect -330 -1550 -250 -1510
rect -330 -1590 -310 -1550
rect -270 -1590 -250 -1550
rect -330 -1630 -250 -1590
rect -330 -1670 -310 -1630
rect -270 -1670 -250 -1630
rect -330 -1710 -250 -1670
rect -330 -1750 -310 -1710
rect -270 -1750 -250 -1710
rect -330 -1790 -250 -1750
rect -330 -1830 -310 -1790
rect -270 -1830 -250 -1790
rect -330 -1850 -250 -1830
rect -150 -1070 -70 -1050
rect -150 -1110 -130 -1070
rect -90 -1110 -70 -1070
rect -150 -1150 -70 -1110
rect -150 -1190 -130 -1150
rect -90 -1190 -70 -1150
rect -150 -1230 -70 -1190
rect -150 -1270 -130 -1230
rect -90 -1270 -70 -1230
rect -150 -1310 -70 -1270
rect -150 -1350 -130 -1310
rect -90 -1350 -70 -1310
rect -150 -1390 -70 -1350
rect -150 -1430 -130 -1390
rect -90 -1430 -70 -1390
rect -150 -1470 -70 -1430
rect -150 -1510 -130 -1470
rect -90 -1510 -70 -1470
rect -150 -1550 -70 -1510
rect -150 -1590 -130 -1550
rect -90 -1590 -70 -1550
rect -150 -1630 -70 -1590
rect -150 -1670 -130 -1630
rect -90 -1670 -70 -1630
rect -150 -1710 -70 -1670
rect -150 -1750 -130 -1710
rect -90 -1750 -70 -1710
rect -150 -1790 -70 -1750
rect -150 -1830 -130 -1790
rect -90 -1830 -70 -1790
rect -150 -1850 -70 -1830
rect 30 -1070 110 -1050
rect 30 -1110 50 -1070
rect 90 -1110 110 -1070
rect 30 -1150 110 -1110
rect 30 -1190 50 -1150
rect 90 -1190 110 -1150
rect 30 -1230 110 -1190
rect 30 -1270 50 -1230
rect 90 -1270 110 -1230
rect 30 -1310 110 -1270
rect 30 -1350 50 -1310
rect 90 -1350 110 -1310
rect 30 -1390 110 -1350
rect 30 -1430 50 -1390
rect 90 -1430 110 -1390
rect 30 -1470 110 -1430
rect 30 -1510 50 -1470
rect 90 -1510 110 -1470
rect 2440 -1080 2520 -1060
rect 2440 -1120 2460 -1080
rect 2500 -1120 2520 -1080
rect 2440 -1160 2520 -1120
rect 2440 -1200 2460 -1160
rect 2500 -1200 2520 -1160
rect 2440 -1240 2520 -1200
rect 2440 -1280 2460 -1240
rect 2500 -1280 2520 -1240
rect 2440 -1320 2520 -1280
rect 2440 -1360 2460 -1320
rect 2500 -1360 2520 -1320
rect 30 -1550 110 -1510
rect 30 -1590 50 -1550
rect 90 -1590 110 -1550
rect 30 -1630 110 -1590
rect 30 -1670 50 -1630
rect 90 -1670 110 -1630
rect 2440 -1400 2520 -1360
rect 2440 -1440 2460 -1400
rect 2500 -1440 2520 -1400
rect 2440 -1480 2520 -1440
rect 2440 -1520 2460 -1480
rect 2500 -1520 2520 -1480
rect 2440 -1560 2520 -1520
rect 2440 -1600 2460 -1560
rect 2500 -1600 2520 -1560
rect 2440 -1640 2520 -1600
rect 30 -1710 110 -1670
rect 30 -1750 50 -1710
rect 90 -1750 110 -1710
rect 30 -1790 110 -1750
rect 30 -1830 50 -1790
rect 90 -1830 110 -1790
rect 30 -1850 110 -1830
rect 2440 -1680 2460 -1640
rect 2500 -1680 2520 -1640
rect 2440 -1720 2520 -1680
rect 2440 -1760 2460 -1720
rect 2500 -1760 2520 -1720
rect 2440 -1800 2520 -1760
rect 2440 -1840 2460 -1800
rect 2500 -1840 2520 -1800
rect 2440 -1860 2520 -1840
rect 2620 -1080 2700 -1060
rect 2620 -1120 2640 -1080
rect 2680 -1120 2700 -1080
rect 2620 -1160 2700 -1120
rect 2620 -1200 2640 -1160
rect 2680 -1200 2700 -1160
rect 2620 -1240 2700 -1200
rect 2620 -1280 2640 -1240
rect 2680 -1280 2700 -1240
rect 2620 -1320 2700 -1280
rect 2620 -1360 2640 -1320
rect 2680 -1360 2700 -1320
rect 2620 -1400 2700 -1360
rect 2620 -1440 2640 -1400
rect 2680 -1440 2700 -1400
rect 2620 -1480 2700 -1440
rect 2620 -1520 2640 -1480
rect 2680 -1520 2700 -1480
rect 2620 -1560 2700 -1520
rect 2620 -1600 2640 -1560
rect 2680 -1600 2700 -1560
rect 2620 -1640 2700 -1600
rect 2620 -1680 2640 -1640
rect 2680 -1680 2700 -1640
rect 2620 -1720 2700 -1680
rect 2620 -1760 2640 -1720
rect 2680 -1760 2700 -1720
rect 2620 -1800 2700 -1760
rect 2620 -1840 2640 -1800
rect 2680 -1840 2700 -1800
rect 2620 -1860 2700 -1840
rect 2800 -1080 2880 -1060
rect 2800 -1120 2820 -1080
rect 2860 -1120 2880 -1080
rect 2800 -1160 2880 -1120
rect 2800 -1200 2820 -1160
rect 2860 -1200 2880 -1160
rect 2800 -1240 2880 -1200
rect 2800 -1280 2820 -1240
rect 2860 -1280 2880 -1240
rect 2800 -1320 2880 -1280
rect 2800 -1360 2820 -1320
rect 2860 -1360 2880 -1320
rect 2800 -1400 2880 -1360
rect 2800 -1440 2820 -1400
rect 2860 -1440 2880 -1400
rect 2800 -1480 2880 -1440
rect 2800 -1520 2820 -1480
rect 2860 -1520 2880 -1480
rect 2800 -1560 2880 -1520
rect 2800 -1600 2820 -1560
rect 2860 -1600 2880 -1560
rect 2800 -1640 2880 -1600
rect 2800 -1680 2820 -1640
rect 2860 -1680 2880 -1640
rect 2800 -1720 2880 -1680
rect 2800 -1760 2820 -1720
rect 2860 -1760 2880 -1720
rect 2800 -1800 2880 -1760
rect 2800 -1840 2820 -1800
rect 2860 -1840 2880 -1800
rect 2800 -1860 2880 -1840
<< ndiffc >>
rect 650 -1150 690 -1110
rect 650 -1230 690 -1190
rect 650 -1310 690 -1270
rect 650 -1390 690 -1350
rect 830 -1150 870 -1110
rect 830 -1230 870 -1190
rect 830 -1310 870 -1270
rect 830 -1390 870 -1350
rect 1010 -1150 1050 -1110
rect 1010 -1230 1050 -1190
rect 1010 -1310 1050 -1270
rect 1010 -1390 1050 -1350
rect 1420 -1210 1460 -1170
rect 1420 -1290 1460 -1250
rect 1420 -1370 1460 -1330
rect 1420 -1450 1460 -1410
rect 1600 -1210 1640 -1170
rect 1600 -1290 1640 -1250
rect 1600 -1370 1640 -1330
rect 1600 -1450 1640 -1410
rect 1780 -1210 1820 -1170
rect 1780 -1290 1820 -1250
rect 1780 -1370 1820 -1330
rect 1780 -1450 1820 -1410
<< pdiffc >>
rect -380 300 -340 340
rect -380 220 -340 260
rect -380 140 -340 180
rect -380 60 -340 100
rect -200 300 -160 340
rect 370 300 410 340
rect -200 220 -160 260
rect -200 140 -160 180
rect -200 60 -160 100
rect 370 220 410 260
rect 370 140 410 180
rect 370 60 410 100
rect 550 300 590 340
rect 550 220 590 260
rect 550 140 590 180
rect 550 60 590 100
rect 730 300 770 340
rect 730 220 770 260
rect 730 140 770 180
rect 730 60 770 100
rect 910 300 950 340
rect 1470 300 1510 340
rect 910 220 950 260
rect 910 140 950 180
rect 910 60 950 100
rect 1470 220 1510 260
rect 1470 140 1510 180
rect 1470 60 1510 100
rect 1650 300 1690 340
rect 1650 220 1690 260
rect 1650 140 1690 180
rect 1650 60 1690 100
rect 1830 300 1870 340
rect 1830 220 1870 260
rect 1830 140 1870 180
rect 1830 60 1870 100
rect 2010 300 2050 340
rect 2570 290 2610 330
rect 2010 220 2050 260
rect 2010 140 2050 180
rect 2010 60 2050 100
rect 2570 210 2610 250
rect 2570 130 2610 170
rect 2570 50 2610 90
rect 2750 290 2790 330
rect 2750 210 2790 250
rect 2750 130 2790 170
rect 2750 50 2790 90
rect -310 -1110 -270 -1070
rect -310 -1190 -270 -1150
rect -310 -1270 -270 -1230
rect -310 -1350 -270 -1310
rect -310 -1430 -270 -1390
rect -310 -1510 -270 -1470
rect -310 -1590 -270 -1550
rect -310 -1670 -270 -1630
rect -310 -1750 -270 -1710
rect -310 -1830 -270 -1790
rect -130 -1110 -90 -1070
rect -130 -1190 -90 -1150
rect -130 -1270 -90 -1230
rect -130 -1350 -90 -1310
rect -130 -1430 -90 -1390
rect -130 -1510 -90 -1470
rect -130 -1590 -90 -1550
rect -130 -1670 -90 -1630
rect -130 -1750 -90 -1710
rect -130 -1830 -90 -1790
rect 50 -1110 90 -1070
rect 50 -1190 90 -1150
rect 50 -1270 90 -1230
rect 50 -1350 90 -1310
rect 50 -1430 90 -1390
rect 50 -1510 90 -1470
rect 2460 -1120 2500 -1080
rect 2460 -1200 2500 -1160
rect 2460 -1280 2500 -1240
rect 2460 -1360 2500 -1320
rect 50 -1590 90 -1550
rect 50 -1670 90 -1630
rect 2460 -1440 2500 -1400
rect 2460 -1520 2500 -1480
rect 2460 -1600 2500 -1560
rect 50 -1750 90 -1710
rect 50 -1830 90 -1790
rect 2460 -1680 2500 -1640
rect 2460 -1760 2500 -1720
rect 2460 -1840 2500 -1800
rect 2640 -1120 2680 -1080
rect 2640 -1200 2680 -1160
rect 2640 -1280 2680 -1240
rect 2640 -1360 2680 -1320
rect 2640 -1440 2680 -1400
rect 2640 -1520 2680 -1480
rect 2640 -1600 2680 -1560
rect 2640 -1680 2680 -1640
rect 2640 -1760 2680 -1720
rect 2640 -1840 2680 -1800
rect 2820 -1120 2860 -1080
rect 2820 -1200 2860 -1160
rect 2820 -1280 2860 -1240
rect 2820 -1360 2860 -1320
rect 2820 -1440 2860 -1400
rect 2820 -1520 2860 -1480
rect 2820 -1600 2860 -1560
rect 2820 -1680 2860 -1640
rect 2820 -1760 2860 -1720
rect 2820 -1840 2860 -1800
<< psubdiff >>
rect 490 -1100 570 -1070
rect 490 -1140 510 -1100
rect 550 -1140 570 -1100
rect 490 -1170 570 -1140
rect 1900 -1420 1980 -1390
rect 1900 -1460 1920 -1420
rect 1960 -1460 1980 -1420
rect 1900 -1490 1980 -1460
rect -1760 -1940 -1660 -1920
rect -1760 -1980 -1730 -1940
rect -1690 -1980 -1660 -1940
rect -1760 -2000 -1660 -1980
<< nsubdiff >>
rect -540 330 -460 360
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect 210 340 290 370
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 1310 270 1390 300
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect 2410 260 2490 290
rect -470 -1070 -390 -1040
rect -470 -1110 -450 -1070
rect -410 -1110 -390 -1070
rect -470 -1140 -390 -1110
rect 2300 -1100 2380 -1070
rect 2300 -1140 2320 -1100
rect 2360 -1140 2380 -1100
rect 2300 -1170 2380 -1140
rect -1480 -1920 -1380 -1900
rect -1480 -1960 -1450 -1920
rect -1410 -1960 -1380 -1920
rect -1480 -1980 -1380 -1960
<< psubdiffcont >>
rect 510 -1140 550 -1100
rect 1920 -1460 1960 -1420
rect -1730 -1980 -1690 -1940
<< nsubdiffcont >>
rect -520 290 -480 330
rect 230 300 270 340
rect 1330 300 1370 340
rect 2430 290 2470 330
rect -450 -1110 -410 -1070
rect 2320 -1140 2360 -1100
rect -1450 -1960 -1410 -1920
<< poly >>
rect -320 510 -220 540
rect -320 470 -270 510
rect -230 470 -220 510
rect -320 360 -220 470
rect 430 510 890 540
rect 430 470 500 510
rect 540 470 600 510
rect 640 470 890 510
rect 430 440 890 470
rect 430 360 530 440
rect 610 360 710 440
rect 790 360 890 440
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 1530 360 1630 440
rect 1710 360 1810 440
rect 1890 360 1990 440
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 350 2730 460
rect -320 -80 -220 0
rect 430 -80 530 0
rect 610 -80 710 0
rect 790 -80 890 0
rect 1530 -80 1630 0
rect 1710 -80 1810 0
rect 1890 -80 1990 0
rect 2630 -90 2730 -10
rect -250 -1050 -150 -970
rect -70 -1050 30 -970
rect 710 -1080 810 -1000
rect 890 -1080 990 -1000
rect 1480 -1080 1580 -1000
rect 1660 -1080 1760 -1000
rect 2520 -1060 2620 -980
rect 2700 -1060 2800 -980
rect 710 -1560 810 -1480
rect 890 -1560 990 -1480
rect 710 -1590 990 -1560
rect 710 -1630 780 -1590
rect 820 -1630 880 -1590
rect 920 -1630 990 -1590
rect 710 -1660 990 -1630
rect 1480 -1560 1580 -1480
rect 1660 -1560 1760 -1480
rect 1480 -1590 1760 -1560
rect 1480 -1630 1560 -1590
rect 1600 -1630 1650 -1590
rect 1690 -1630 1760 -1590
rect 1480 -1660 1760 -1630
rect -250 -1930 -150 -1850
rect -70 -1930 30 -1850
rect -250 -1960 30 -1930
rect -250 -2000 -240 -1960
rect -200 -2000 -20 -1960
rect 20 -2000 30 -1960
rect -250 -2030 30 -2000
rect 2520 -1940 2620 -1860
rect 2700 -1940 2800 -1860
rect 2520 -1970 2800 -1940
rect 2520 -2010 2530 -1970
rect 2570 -2010 2750 -1970
rect 2790 -2010 2800 -1970
rect 2520 -2040 2800 -2010
<< polycont >>
rect -270 470 -230 510
rect 500 470 540 510
rect 600 470 640 510
rect 1560 470 1600 510
rect 1740 470 1780 510
rect 1920 470 1960 510
rect 2660 460 2700 500
rect 780 -1630 820 -1590
rect 880 -1630 920 -1590
rect 1560 -1630 1600 -1590
rect 1650 -1630 1690 -1590
rect -240 -2000 -200 -1960
rect -20 -2000 20 -1960
rect 2530 -2010 2570 -1970
rect 2750 -2010 2790 -1970
<< locali >>
rect -540 730 790 740
rect -540 680 -520 730
rect -470 680 -390 730
rect -340 680 790 730
rect -540 660 790 680
rect -540 330 -460 660
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect -400 340 -320 660
rect -280 510 -220 540
rect -280 470 -270 510
rect -230 470 -220 510
rect -280 440 -220 470
rect -400 300 -380 340
rect -340 300 -320 340
rect -400 260 -320 300
rect -400 220 -380 260
rect -340 220 -320 260
rect -400 180 -320 220
rect -400 140 -380 180
rect -340 140 -320 180
rect -400 100 -320 140
rect -400 60 -380 100
rect -340 60 -320 100
rect -400 0 -320 60
rect -220 340 -140 360
rect -220 300 -200 340
rect -160 300 -140 340
rect -220 260 -140 300
rect 210 340 290 660
rect 470 510 670 540
rect 470 470 500 510
rect 540 470 600 510
rect 640 470 670 510
rect 470 440 670 470
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 350 340 430 360
rect 350 300 370 340
rect 410 300 430 340
rect -220 220 -200 260
rect -160 220 -140 260
rect -220 180 -140 220
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 0 -140 60
rect 350 260 430 300
rect 350 220 370 260
rect 410 220 430 260
rect 350 180 430 220
rect 350 140 370 180
rect 410 140 430 180
rect 350 100 430 140
rect 350 60 370 100
rect 410 60 430 100
rect 350 0 430 60
rect 530 340 610 360
rect 530 300 550 340
rect 590 300 610 340
rect 530 260 610 300
rect 530 220 550 260
rect 590 220 610 260
rect 530 180 610 220
rect 530 140 550 180
rect 590 140 610 180
rect 530 100 610 140
rect 530 60 550 100
rect 590 60 610 100
rect 530 0 610 60
rect 710 340 790 660
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 430 2730 460
rect 710 300 730 340
rect 770 300 790 340
rect 710 260 790 300
rect 710 220 730 260
rect 770 220 790 260
rect 710 180 790 220
rect 710 140 730 180
rect 770 140 790 180
rect 710 100 790 140
rect 710 60 730 100
rect 770 60 790 100
rect 710 0 790 60
rect 890 340 970 360
rect 890 300 910 340
rect 950 300 970 340
rect 890 260 970 300
rect 890 220 910 260
rect 950 220 970 260
rect 890 180 970 220
rect 890 140 910 180
rect 950 140 970 180
rect 890 100 970 140
rect 890 60 910 100
rect 950 60 970 100
rect 890 -150 970 60
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 1310 -150 1390 300
rect 1450 340 1530 360
rect 1450 300 1470 340
rect 1510 300 1530 340
rect 1450 260 1530 300
rect 1450 220 1470 260
rect 1510 220 1530 260
rect 1450 180 1530 220
rect 1450 140 1470 180
rect 1510 140 1530 180
rect 1450 100 1530 140
rect 1450 60 1470 100
rect 1510 60 1530 100
rect 1450 -150 1530 60
rect 890 -230 1530 -150
rect 1630 340 1710 360
rect 1630 300 1650 340
rect 1690 300 1710 340
rect 1630 260 1710 300
rect 1630 220 1650 260
rect 1690 220 1710 260
rect 1630 180 1710 220
rect 1630 140 1650 180
rect 1690 140 1710 180
rect 1630 100 1710 140
rect 1630 60 1650 100
rect 1690 60 1710 100
rect 1630 -540 1710 60
rect 1810 340 1890 360
rect 1810 300 1830 340
rect 1870 300 1890 340
rect 1810 260 1890 300
rect 1810 220 1830 260
rect 1870 220 1890 260
rect 1810 180 1890 220
rect 1810 140 1830 180
rect 1870 140 1890 180
rect 1810 100 1890 140
rect 1810 60 1830 100
rect 1870 60 1890 100
rect 1810 0 1890 60
rect 1990 340 2070 360
rect 1990 300 2010 340
rect 2050 300 2070 340
rect 1990 260 2070 300
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect 2410 260 2490 290
rect 2550 330 2630 350
rect 2550 290 2570 330
rect 2610 290 2630 330
rect 1990 220 2010 260
rect 2050 220 2070 260
rect 1990 180 2070 220
rect 1990 140 2010 180
rect 2050 140 2070 180
rect 1990 100 2070 140
rect 1990 60 2010 100
rect 2050 60 2070 100
rect 1990 0 2070 60
rect 2550 250 2630 290
rect 2550 210 2570 250
rect 2610 210 2630 250
rect 2550 170 2630 210
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -10 2630 50
rect 2730 330 2810 350
rect 2730 290 2750 330
rect 2790 290 2810 330
rect 2730 250 2810 290
rect 2730 210 2750 250
rect 2790 210 2810 250
rect 2730 170 2810 210
rect 2730 130 2750 170
rect 2790 130 2810 170
rect 2730 90 2810 130
rect 2730 50 2750 90
rect 2790 50 3220 90
rect 2730 -10 3220 50
rect 10 -640 2380 -540
rect 10 -740 110 -640
rect -470 -840 110 -740
rect -470 -1070 -390 -840
rect -470 -1110 -450 -1070
rect -410 -1110 -390 -1070
rect -470 -1140 -390 -1110
rect -330 -1070 -250 -1050
rect -330 -1110 -310 -1070
rect -270 -1110 -250 -1070
rect -330 -1150 -250 -1110
rect -330 -1190 -310 -1150
rect -270 -1190 -250 -1150
rect -330 -1230 -250 -1190
rect -330 -1270 -310 -1230
rect -270 -1270 -250 -1230
rect -330 -1310 -250 -1270
rect -330 -1350 -310 -1310
rect -270 -1350 -250 -1310
rect -330 -1390 -250 -1350
rect -330 -1430 -310 -1390
rect -270 -1430 -250 -1390
rect -330 -1470 -250 -1430
rect -330 -1510 -310 -1470
rect -270 -1510 -250 -1470
rect -330 -1550 -250 -1510
rect -330 -1590 -310 -1550
rect -270 -1590 -250 -1550
rect -330 -1630 -250 -1590
rect -330 -1670 -310 -1630
rect -270 -1670 -250 -1630
rect -330 -1710 -250 -1670
rect -1760 -1940 -1660 -1920
rect -1760 -1980 -1730 -1940
rect -1690 -1980 -1660 -1940
rect -1760 -2000 -1660 -1980
rect -1590 -2020 -1550 -1720
rect -330 -1750 -310 -1710
rect -270 -1750 -250 -1710
rect -330 -1790 -250 -1750
rect -330 -1830 -310 -1790
rect -270 -1830 -250 -1790
rect -330 -1850 -250 -1830
rect -150 -1070 -70 -1050
rect -150 -1110 -130 -1070
rect -90 -1110 -70 -1070
rect -150 -1150 -70 -1110
rect -150 -1190 -130 -1150
rect -90 -1190 -70 -1150
rect -150 -1230 -70 -1190
rect -150 -1270 -130 -1230
rect -90 -1270 -70 -1230
rect -150 -1310 -70 -1270
rect -150 -1350 -130 -1310
rect -90 -1350 -70 -1310
rect -150 -1390 -70 -1350
rect -150 -1430 -130 -1390
rect -90 -1430 -70 -1390
rect -150 -1470 -70 -1430
rect -150 -1510 -130 -1470
rect -90 -1510 -70 -1470
rect -150 -1550 -70 -1510
rect -150 -1590 -130 -1550
rect -90 -1590 -70 -1550
rect -150 -1630 -70 -1590
rect -150 -1670 -130 -1630
rect -90 -1670 -70 -1630
rect -150 -1710 -70 -1670
rect -150 -1750 -130 -1710
rect -90 -1750 -70 -1710
rect -150 -1790 -70 -1750
rect -150 -1830 -130 -1790
rect -90 -1830 -70 -1790
rect -1480 -1920 -1380 -1900
rect -1480 -1960 -1450 -1920
rect -1410 -1960 -1380 -1920
rect -250 -1940 -190 -1930
rect -1480 -1980 -1380 -1960
rect -1110 -1960 -190 -1940
rect -1110 -2000 -240 -1960
rect -200 -2000 -190 -1960
rect -1110 -2020 -190 -2000
rect -1590 -2100 -1030 -2020
rect -250 -2030 -190 -2020
rect -1590 -2180 -1550 -2100
rect -150 -2170 -70 -1830
rect 30 -1070 110 -840
rect 30 -1110 50 -1070
rect 90 -1110 110 -1070
rect 30 -1150 110 -1110
rect 30 -1190 50 -1150
rect 90 -1190 110 -1150
rect 490 -1100 570 -1070
rect 490 -1140 510 -1100
rect 550 -1140 570 -1100
rect 490 -1170 570 -1140
rect 630 -1110 710 -1080
rect 630 -1150 650 -1110
rect 690 -1150 710 -1110
rect 30 -1230 110 -1190
rect 30 -1270 50 -1230
rect 90 -1270 110 -1230
rect 30 -1310 110 -1270
rect 30 -1350 50 -1310
rect 90 -1350 110 -1310
rect 30 -1390 110 -1350
rect 30 -1430 50 -1390
rect 90 -1430 110 -1390
rect 30 -1470 110 -1430
rect 30 -1510 50 -1470
rect 90 -1510 110 -1470
rect 30 -1550 110 -1510
rect 30 -1590 50 -1550
rect 90 -1590 110 -1550
rect 30 -1630 110 -1590
rect 30 -1670 50 -1630
rect 90 -1670 110 -1630
rect 30 -1710 110 -1670
rect 30 -1750 50 -1710
rect 90 -1750 110 -1710
rect 30 -1790 110 -1750
rect 30 -1830 50 -1790
rect 90 -1830 110 -1790
rect 30 -1850 110 -1830
rect 630 -1190 710 -1150
rect 630 -1230 650 -1190
rect 690 -1230 710 -1190
rect 630 -1270 710 -1230
rect 630 -1310 650 -1270
rect 690 -1310 710 -1270
rect 630 -1350 710 -1310
rect 630 -1390 650 -1350
rect 690 -1390 710 -1350
rect -30 -1960 30 -1930
rect -30 -2000 -20 -1960
rect 20 -2000 30 -1960
rect -30 -2030 30 -2000
rect 630 -2170 710 -1390
rect 810 -1110 890 -640
rect 810 -1150 830 -1110
rect 870 -1150 890 -1110
rect 810 -1190 890 -1150
rect 810 -1230 830 -1190
rect 870 -1230 890 -1190
rect 810 -1270 890 -1230
rect 810 -1310 830 -1270
rect 870 -1310 890 -1270
rect 810 -1350 890 -1310
rect 810 -1390 830 -1350
rect 870 -1390 890 -1350
rect 810 -1480 890 -1390
rect 990 -1110 1070 -1080
rect 990 -1150 1010 -1110
rect 1050 -1150 1070 -1110
rect 990 -1190 1070 -1150
rect 990 -1230 1010 -1190
rect 1050 -1230 1070 -1190
rect 990 -1270 1070 -1230
rect 990 -1310 1010 -1270
rect 1050 -1310 1070 -1270
rect 990 -1350 1070 -1310
rect 990 -1390 1010 -1350
rect 1050 -1390 1070 -1350
rect 990 -1480 1070 -1390
rect 1400 -1170 1480 -1080
rect 1400 -1210 1420 -1170
rect 1460 -1210 1480 -1170
rect 1400 -1250 1480 -1210
rect 1400 -1290 1420 -1250
rect 1460 -1290 1480 -1250
rect 1400 -1330 1480 -1290
rect 1400 -1370 1420 -1330
rect 1460 -1370 1480 -1330
rect 1400 -1410 1480 -1370
rect 1400 -1450 1420 -1410
rect 1460 -1450 1480 -1410
rect 1400 -1480 1480 -1450
rect 1580 -1170 1660 -640
rect 2300 -740 2380 -640
rect 2300 -840 2520 -740
rect 1580 -1210 1600 -1170
rect 1640 -1210 1660 -1170
rect 1580 -1250 1660 -1210
rect 1580 -1290 1600 -1250
rect 1640 -1290 1660 -1250
rect 1580 -1330 1660 -1290
rect 1580 -1370 1600 -1330
rect 1640 -1370 1660 -1330
rect 1580 -1410 1660 -1370
rect 1580 -1450 1600 -1410
rect 1640 -1450 1660 -1410
rect 1580 -1480 1660 -1450
rect 1760 -1170 1840 -1080
rect 2300 -1100 2380 -840
rect 2300 -1140 2320 -1100
rect 2360 -1140 2380 -1100
rect 2300 -1170 2380 -1140
rect 2440 -1080 2520 -840
rect 2440 -1120 2460 -1080
rect 2500 -1120 2520 -1080
rect 2440 -1160 2520 -1120
rect 1760 -1210 1780 -1170
rect 1820 -1210 1840 -1170
rect 1760 -1250 1840 -1210
rect 1760 -1290 1780 -1250
rect 1820 -1290 1840 -1250
rect 1760 -1330 1840 -1290
rect 1760 -1370 1780 -1330
rect 1820 -1370 1840 -1330
rect 1760 -1410 1840 -1370
rect 2440 -1200 2460 -1160
rect 2500 -1200 2520 -1160
rect 2440 -1240 2520 -1200
rect 2440 -1280 2460 -1240
rect 2500 -1280 2520 -1240
rect 2440 -1320 2520 -1280
rect 2440 -1360 2460 -1320
rect 2500 -1360 2520 -1320
rect 1760 -1450 1780 -1410
rect 1820 -1450 1840 -1410
rect 750 -1590 950 -1560
rect 750 -1630 780 -1590
rect 820 -1630 880 -1590
rect 920 -1630 950 -1590
rect 750 -1660 950 -1630
rect 1540 -1590 1710 -1560
rect 1540 -1630 1560 -1590
rect 1600 -1630 1650 -1590
rect 1690 -1630 1710 -1590
rect 1540 -1660 1710 -1630
rect -150 -2190 710 -2170
rect -150 -2230 -130 -2190
rect -90 -2230 710 -2190
rect -150 -2250 710 -2230
rect 810 -2330 890 -1660
rect 1760 -2100 1840 -1450
rect 1900 -1420 1980 -1390
rect 1900 -1460 1920 -1420
rect 1960 -1460 1980 -1420
rect 1900 -1490 1980 -1460
rect 2440 -1400 2520 -1360
rect 2440 -1440 2460 -1400
rect 2500 -1440 2520 -1400
rect 2440 -1480 2520 -1440
rect 2440 -1520 2460 -1480
rect 2500 -1520 2520 -1480
rect 2440 -1560 2520 -1520
rect 2440 -1600 2460 -1560
rect 2500 -1600 2520 -1560
rect 2440 -1640 2520 -1600
rect 2440 -1680 2460 -1640
rect 2500 -1680 2520 -1640
rect 2440 -1720 2520 -1680
rect 2440 -1760 2460 -1720
rect 2500 -1760 2520 -1720
rect 2440 -1800 2520 -1760
rect 2440 -1840 2460 -1800
rect 2500 -1840 2520 -1800
rect 2440 -1860 2520 -1840
rect 2620 -1080 2700 -1060
rect 2620 -1120 2640 -1080
rect 2680 -1120 2700 -1080
rect 2620 -1160 2700 -1120
rect 2620 -1200 2640 -1160
rect 2680 -1200 2700 -1160
rect 2620 -1240 2700 -1200
rect 2620 -1280 2640 -1240
rect 2680 -1280 2700 -1240
rect 2620 -1320 2700 -1280
rect 2620 -1360 2640 -1320
rect 2680 -1360 2700 -1320
rect 2620 -1400 2700 -1360
rect 2620 -1440 2640 -1400
rect 2680 -1440 2700 -1400
rect 2620 -1480 2700 -1440
rect 2620 -1520 2640 -1480
rect 2680 -1520 2700 -1480
rect 2620 -1560 2700 -1520
rect 2620 -1600 2640 -1560
rect 2680 -1600 2700 -1560
rect 2620 -1640 2700 -1600
rect 2620 -1680 2640 -1640
rect 2680 -1680 2700 -1640
rect 2620 -1720 2700 -1680
rect 2620 -1760 2640 -1720
rect 2680 -1760 2700 -1720
rect 2620 -1800 2700 -1760
rect 2620 -1840 2640 -1800
rect 2680 -1840 2700 -1800
rect 2520 -1970 2580 -1940
rect 2520 -2010 2530 -1970
rect 2570 -2010 2580 -1970
rect 2520 -2040 2580 -2010
rect 2620 -2100 2700 -1840
rect 2800 -1080 2880 -1060
rect 2800 -1120 2820 -1080
rect 2860 -1120 2880 -1080
rect 2800 -1160 2880 -1120
rect 2800 -1200 2820 -1160
rect 2860 -1200 2880 -1160
rect 2800 -1240 2880 -1200
rect 2800 -1280 2820 -1240
rect 2860 -1280 2880 -1240
rect 2800 -1320 2880 -1280
rect 2800 -1360 2820 -1320
rect 2860 -1360 2880 -1320
rect 2800 -1400 2880 -1360
rect 2800 -1440 2820 -1400
rect 2860 -1440 2880 -1400
rect 2800 -1480 2880 -1440
rect 2800 -1520 2820 -1480
rect 2860 -1520 2880 -1480
rect 2800 -1560 2880 -1520
rect 2800 -1600 2820 -1560
rect 2860 -1600 2880 -1560
rect 2800 -1640 2880 -1600
rect 2800 -1680 2820 -1640
rect 2860 -1680 2880 -1640
rect 2800 -1720 2880 -1680
rect 2800 -1760 2820 -1720
rect 2860 -1760 2880 -1720
rect 2800 -1800 2880 -1760
rect 2800 -1840 2820 -1800
rect 2860 -1840 2880 -1800
rect 2800 -1860 2880 -1840
rect 2740 -1970 2800 -1940
rect 2740 -2010 2750 -1970
rect 2790 -2010 2800 -1970
rect 2740 -2040 2800 -2010
rect 3120 -2100 3220 -10
rect 1760 -2200 3220 -2100
rect -1110 -2360 2880 -2330
rect -1110 -2400 2820 -2360
rect 2860 -2400 2880 -2360
rect -1110 -2430 2880 -2400
rect -1110 -2550 -1010 -2430
rect -1540 -2580 -1010 -2550
rect -1540 -2620 -1510 -2580
rect -1470 -2620 -1010 -2580
rect -1540 -2650 -1010 -2620
rect -400 -2600 570 -2580
rect -400 -2640 -380 -2600
rect -340 -2640 510 -2600
rect 550 -2640 570 -2600
rect -400 -2660 570 -2640
rect -40 -3080 40 -3060
rect -40 -3120 -20 -3080
rect 20 -3120 40 -3080
rect 2510 -3090 2690 -2920
rect 2630 -3120 2690 -3090
rect -40 -3140 40 -3120
<< viali >>
rect -520 680 -470 730
rect -390 680 -340 730
rect -520 290 -480 330
rect -270 470 -230 510
rect 500 470 540 510
rect 600 470 640 510
rect 230 300 270 340
rect 370 300 410 340
rect -200 140 -160 180
rect -200 60 -160 100
rect 370 220 410 260
rect 550 60 590 100
rect 1560 470 1600 510
rect 1740 470 1780 510
rect 1920 470 1960 510
rect 2660 460 2700 500
rect 730 300 770 340
rect 730 220 770 260
rect 910 60 950 100
rect 1330 300 1370 340
rect 1470 300 1510 340
rect 1470 220 1510 260
rect 1650 60 1690 100
rect 1830 300 1870 340
rect 1830 220 1870 260
rect 2430 290 2470 330
rect 2010 60 2050 100
rect 2570 130 2610 170
rect 2570 50 2610 90
rect -450 -1110 -410 -1070
rect -310 -1110 -270 -1070
rect -310 -1190 -270 -1150
rect -1600 -1560 -1560 -1520
rect -1730 -1980 -1690 -1940
rect -310 -1750 -270 -1710
rect -310 -1830 -270 -1790
rect -1450 -1960 -1410 -1920
rect -240 -2000 -200 -1960
rect 50 -1110 90 -1070
rect 50 -1190 90 -1150
rect 510 -1140 550 -1100
rect 650 -1150 690 -1110
rect 50 -1750 90 -1710
rect 50 -1830 90 -1790
rect 650 -1230 690 -1190
rect -20 -2000 20 -1960
rect 1010 -1150 1050 -1110
rect 1010 -1230 1050 -1190
rect 1420 -1210 1460 -1170
rect 1420 -1290 1460 -1250
rect 2320 -1140 2360 -1100
rect 2460 -1120 2500 -1080
rect 1780 -1210 1820 -1170
rect 1780 -1290 1820 -1250
rect 2460 -1200 2500 -1160
rect 780 -1630 820 -1590
rect 880 -1630 920 -1590
rect 1560 -1630 1600 -1590
rect 1650 -1630 1690 -1590
rect -130 -2230 -90 -2190
rect -1510 -2310 -1470 -2270
rect -1430 -2310 -1390 -2270
rect 1920 -1460 1960 -1420
rect 2460 -1760 2500 -1720
rect 2460 -1840 2500 -1800
rect 2530 -2010 2570 -1970
rect 2820 -1120 2860 -1080
rect 2820 -1200 2860 -1160
rect 2820 -1760 2860 -1720
rect 2820 -1840 2860 -1800
rect 2750 -2010 2790 -1970
rect 2820 -2400 2860 -2360
rect -1510 -2620 -1470 -2580
rect -380 -2640 -340 -2600
rect 510 -2640 550 -2600
rect -20 -3120 20 -3080
<< metal1 >>
rect -1320 730 -320 740
rect -1320 680 -520 730
rect -470 680 -390 730
rect -340 680 -320 730
rect -1320 660 -320 680
rect -1620 -1520 -1540 -1340
rect -1320 -1490 -1220 660
rect -320 510 -220 540
rect -320 470 -270 510
rect -230 470 -220 510
rect -320 440 -220 470
rect 430 510 890 540
rect 430 470 500 510
rect 540 470 600 510
rect 640 470 890 510
rect 430 440 890 470
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 430 2730 460
rect -540 330 -460 360
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect 210 340 290 370
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 350 340 430 360
rect 350 300 370 340
rect 410 330 430 340
rect 710 340 790 360
rect 710 330 730 340
rect 410 300 730 330
rect 770 300 790 340
rect 350 260 790 300
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 1310 270 1390 300
rect 1450 340 1530 360
rect 1810 340 1890 360
rect 1450 300 1470 340
rect 1510 300 1830 340
rect 1870 300 1890 340
rect 350 220 370 260
rect 410 230 730 260
rect 410 220 430 230
rect 350 200 430 220
rect 710 220 730 230
rect 770 220 790 260
rect 710 200 790 220
rect 1450 260 1890 300
rect 1450 220 1470 260
rect 1510 230 1830 260
rect 1510 220 1530 230
rect 1450 200 1530 220
rect 1810 220 1830 230
rect 1870 220 1890 260
rect 1810 200 1890 220
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect -220 180 -140 200
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 -380 -140 60
rect 530 100 970 120
rect 530 60 550 100
rect 590 60 910 100
rect 950 60 970 100
rect 530 20 970 60
rect 530 0 610 20
rect 890 0 970 20
rect 1630 100 2070 120
rect 1630 60 1650 100
rect 1690 60 2010 100
rect 2050 60 2070 100
rect 1630 0 2070 60
rect 2410 -380 2490 290
rect 2550 170 2630 190
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -380 2630 50
rect -220 -460 2630 -380
rect 230 -930 1310 -830
rect -470 -1070 -390 -1040
rect -470 -1110 -450 -1070
rect -410 -1110 -390 -1070
rect -470 -1140 -390 -1110
rect -330 -1070 -250 -1050
rect -330 -1110 -310 -1070
rect -270 -1080 -250 -1070
rect 30 -1070 110 -1050
rect 30 -1080 50 -1070
rect -270 -1110 50 -1080
rect 90 -1110 110 -1070
rect -330 -1150 110 -1110
rect -330 -1190 -310 -1150
rect -270 -1180 50 -1150
rect -270 -1190 -250 -1180
rect -330 -1210 -250 -1190
rect 30 -1190 50 -1180
rect 90 -1190 110 -1150
rect 30 -1210 110 -1190
rect -1620 -1560 -1600 -1520
rect -1560 -1560 -1540 -1520
rect -1620 -1580 -1540 -1560
rect -330 -1710 -250 -1690
rect -330 -1750 -310 -1710
rect -270 -1720 -250 -1710
rect 30 -1710 110 -1690
rect 30 -1720 50 -1710
rect -270 -1750 50 -1720
rect 90 -1750 110 -1710
rect -330 -1790 110 -1750
rect -330 -1830 -310 -1790
rect -270 -1820 50 -1790
rect -270 -1830 -250 -1820
rect -330 -1850 -250 -1830
rect 30 -1830 50 -1820
rect 90 -1830 110 -1790
rect 30 -1850 110 -1830
rect -1860 -1920 -1760 -1850
rect -1320 -1900 -1220 -1850
rect -1480 -1920 -1220 -1900
rect -1860 -1940 -1660 -1920
rect -1860 -1980 -1730 -1940
rect -1690 -1980 -1660 -1940
rect -1480 -1960 -1450 -1920
rect -1410 -1960 -1220 -1920
rect 230 -1930 330 -930
rect -1480 -1980 -1220 -1960
rect -1860 -2000 -1660 -1980
rect -1860 -2150 -1760 -2000
rect -1320 -2150 -1220 -1980
rect -250 -1960 330 -1930
rect -250 -2000 -240 -1960
rect -200 -2000 -20 -1960
rect 20 -2000 330 -1960
rect -250 -2030 330 -2000
rect 490 -1100 570 -1070
rect 490 -1140 510 -1100
rect 550 -1140 570 -1100
rect 490 -1870 570 -1140
rect 630 -1110 710 -1080
rect 630 -1150 650 -1110
rect 690 -1120 710 -1110
rect 990 -1110 1070 -1080
rect 990 -1120 1010 -1110
rect 690 -1150 1010 -1120
rect 1050 -1150 1070 -1110
rect 630 -1190 1070 -1150
rect 630 -1230 650 -1190
rect 690 -1220 1010 -1190
rect 690 -1230 710 -1220
rect 630 -1250 710 -1230
rect 990 -1230 1010 -1220
rect 1050 -1230 1070 -1190
rect 990 -1250 1070 -1230
rect 1210 -1560 1310 -930
rect 1400 -1170 1480 -1080
rect 1400 -1210 1420 -1170
rect 1460 -1180 1480 -1170
rect 1760 -1170 1840 -1080
rect 2300 -1100 2380 -1070
rect 2300 -1140 2320 -1100
rect 2360 -1140 2380 -1100
rect 2300 -1170 2380 -1140
rect 2440 -1080 2520 -1060
rect 2440 -1120 2460 -1080
rect 2500 -1090 2520 -1080
rect 2800 -1080 2880 -1060
rect 2800 -1090 2820 -1080
rect 2500 -1120 2820 -1090
rect 2860 -1120 2880 -1080
rect 2440 -1160 2880 -1120
rect 1760 -1180 1780 -1170
rect 1460 -1210 1780 -1180
rect 1820 -1210 1840 -1170
rect 1400 -1250 1840 -1210
rect 2440 -1200 2460 -1160
rect 2500 -1190 2820 -1160
rect 2500 -1200 2520 -1190
rect 2440 -1220 2520 -1200
rect 2800 -1200 2820 -1190
rect 2860 -1200 2880 -1160
rect 2800 -1220 2880 -1200
rect 1400 -1290 1420 -1250
rect 1460 -1280 1780 -1250
rect 1460 -1290 1480 -1280
rect 1400 -1310 1480 -1290
rect 1760 -1290 1780 -1280
rect 1820 -1290 1840 -1250
rect 1760 -1310 1840 -1290
rect 1900 -1420 1980 -1390
rect 1900 -1460 1920 -1420
rect 1960 -1460 1980 -1420
rect 710 -1590 990 -1560
rect 710 -1630 780 -1590
rect 820 -1630 880 -1590
rect 920 -1630 990 -1590
rect 710 -1660 990 -1630
rect 1210 -1590 1760 -1560
rect 1210 -1630 1560 -1590
rect 1600 -1630 1650 -1590
rect 1690 -1630 1760 -1590
rect 1210 -1660 1760 -1630
rect 1900 -1870 1980 -1460
rect 2440 -1720 2520 -1700
rect 2440 -1760 2460 -1720
rect 2500 -1730 2520 -1720
rect 2800 -1720 2880 -1700
rect 2800 -1730 2820 -1720
rect 2500 -1760 2820 -1730
rect 2860 -1760 2880 -1720
rect 2440 -1800 2880 -1760
rect 2440 -1840 2460 -1800
rect 2500 -1830 2820 -1800
rect 2500 -1840 2520 -1830
rect 2440 -1860 2520 -1840
rect 2800 -1840 2820 -1830
rect 2860 -1840 2880 -1800
rect 2800 -1860 2880 -1840
rect 490 -1950 1980 -1870
rect -190 -2190 -30 -2140
rect -190 -2230 -130 -2190
rect -90 -2230 -30 -2190
rect -1540 -2270 -1370 -2250
rect -1540 -2310 -1510 -2270
rect -1470 -2310 -1430 -2270
rect -1390 -2310 -1370 -2270
rect -190 -2280 -30 -2230
rect -1540 -2320 -1370 -2310
rect -1850 -3060 -1770 -2390
rect -1540 -2580 -1440 -2320
rect -1540 -2620 -1510 -2580
rect -1470 -2620 -1440 -2580
rect -1540 -2650 -1440 -2620
rect -400 -2600 -320 -2580
rect -400 -2640 -380 -2600
rect -340 -2640 -320 -2600
rect -400 -3060 -320 -2640
rect -150 -2920 -70 -2280
rect 490 -2600 570 -1950
rect 2520 -1970 2880 -1940
rect 2520 -2010 2530 -1970
rect 2570 -2010 2750 -1970
rect 2790 -2010 2880 -1970
rect 2520 -2040 2880 -2010
rect 2800 -2360 2880 -2040
rect 2800 -2400 2820 -2360
rect 2860 -2400 2880 -2360
rect 2800 -2430 2880 -2400
rect 490 -2640 510 -2600
rect 550 -2640 570 -2600
rect 490 -2660 570 -2640
rect -150 -3000 350 -2920
rect -1850 -3080 40 -3060
rect -1850 -3120 -20 -3080
rect 20 -3120 40 -3080
rect -1850 -3140 40 -3120
use sky130_fd_pr__res_xhigh_po_0p35_RSCMUS  sky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0
timestamp 1726720190
transform 0 -1 1378 1 0 -2959
box -201 -1438 201 1438
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -1812 -1 0 -1488
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -1812 -1 0 -2148
box -38 -48 314 592
<< labels >>
rlabel metal1 -240 540 -240 540 1 Vbs1
port 1 n
rlabel metal1 2680 530 2680 530 1 Vbs2
port 2 n
rlabel metal1 570 540 570 540 1 Vbs3
port 3 n
rlabel metal1 1770 540 1770 540 1 Vbs4
port 4 n
rlabel metal1 -1540 -1370 -1540 -1370 3 Dctrl
port 5 e
rlabel locali 3060 -2100 3060 -2100 1 Isup
port 6 n
rlabel metal1 -1250 740 -1250 740 1 VDDA
port 7 n
rlabel metal1 -360 -2580 -360 -2580 1 GND
port 8 n
<< end >>
