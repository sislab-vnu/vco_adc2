magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -860 -780 2690 -440
rect -850 -1500 -670 -1480
rect -850 -1810 -690 -1500
rect -850 -1820 -680 -1810
rect 1610 -1910 1810 -1580
rect -190 -2840 -20 -2820
rect 1960 -2830 2320 -2820
rect -190 -3140 -40 -2840
rect 1960 -3140 2280 -2830
rect -190 -3150 -20 -3140
rect 1960 -3150 2350 -3140
<< pwell >>
rect -846 -1006 -714 -854
rect -836 -2046 -704 -1894
rect 1634 -2146 1786 -2014
rect 2114 -2716 2266 -2584
<< psubdiff >>
rect -820 -913 -740 -880
rect -820 -947 -797 -913
rect -763 -947 -740 -913
rect -820 -980 -740 -947
rect -810 -1953 -730 -1920
rect -810 -1987 -787 -1953
rect -753 -1987 -730 -1953
rect -810 -2020 -730 -1987
rect 1660 -2063 1760 -2040
rect 1660 -2097 1693 -2063
rect 1727 -2097 1760 -2063
rect 1660 -2120 1760 -2097
rect 2140 -2633 2240 -2610
rect 2140 -2667 2173 -2633
rect 2207 -2667 2240 -2633
rect 2140 -2690 2240 -2667
<< nsubdiff >>
rect -210 -593 -130 -560
rect -210 -627 -187 -593
rect -153 -627 -130 -593
rect -210 -660 -130 -627
rect -810 -1603 -730 -1570
rect -810 -1637 -787 -1603
rect -753 -1637 -730 -1603
rect -810 -1670 -730 -1637
rect 1680 -1753 1760 -1720
rect 1680 -1787 1703 -1753
rect 1737 -1787 1760 -1753
rect 1680 -1820 1760 -1787
rect -130 -2943 -50 -2910
rect -130 -2977 -107 -2943
rect -73 -2977 -50 -2943
rect -130 -3010 -50 -2977
<< psubdiffcont >>
rect -797 -947 -763 -913
rect -787 -1987 -753 -1953
rect 1693 -2097 1727 -2063
rect 2173 -2667 2207 -2633
<< nsubdiffcont >>
rect -187 -627 -153 -593
rect -787 -1637 -753 -1603
rect 1703 -1787 1737 -1753
rect -107 -2977 -73 -2943
<< locali >>
rect 2630 -540 3140 -470
rect -210 -593 -130 -560
rect -210 -627 -187 -593
rect -153 -627 -130 -593
rect -210 -660 -130 -627
rect 360 -753 400 -750
rect -880 -830 -610 -760
rect -440 -810 20 -770
rect 360 -787 363 -753
rect 397 -787 400 -753
rect 360 -790 400 -787
rect 1820 -783 2300 -760
rect 1820 -817 2103 -783
rect 2137 -817 2300 -783
rect 1820 -840 2300 -817
rect -820 -913 -740 -880
rect -820 -947 -797 -913
rect -763 -947 -740 -913
rect -820 -980 -740 -947
rect -360 -1080 -10 -980
rect 1910 -1080 2280 -990
rect -810 -1603 -730 -1570
rect -430 -1580 1000 -1510
rect -810 -1637 -787 -1603
rect -753 -1637 -730 -1603
rect 930 -1620 1000 -1580
rect 3070 -1610 3140 -540
rect -810 -1670 -730 -1637
rect 2190 -1680 3140 -1610
rect 1680 -1753 1760 -1720
rect 1680 -1787 1703 -1753
rect 1737 -1787 1760 -1753
rect -638 -1817 -598 -1814
rect -638 -1851 -635 -1817
rect -601 -1851 -598 -1817
rect 1680 -1820 1760 -1787
rect 2064 -1773 2104 -1770
rect 2064 -1807 2067 -1773
rect 2101 -1807 2104 -1773
rect 2064 -1810 2104 -1807
rect -638 -1854 -598 -1851
rect 1460 -1900 1800 -1890
rect -810 -1953 -730 -1920
rect 1460 -1940 1870 -1900
rect 2090 -1950 2100 -1940
rect -810 -1987 -787 -1953
rect -753 -1987 -730 -1953
rect -810 -2020 -730 -1987
rect -430 -2033 510 -2020
rect -430 -2067 453 -2033
rect 487 -2067 510 -2033
rect -430 -2090 510 -2067
rect 440 -2130 510 -2090
rect 1660 -2063 1760 -2040
rect 1660 -2097 1693 -2063
rect 1727 -2097 1760 -2063
rect 1660 -2120 1760 -2097
rect 440 -2200 970 -2130
rect -250 -2610 10 -2520
rect 440 -2565 510 -2200
rect 1920 -2610 2350 -2540
rect 2140 -2633 2240 -2610
rect 2140 -2667 2173 -2633
rect 2207 -2667 2240 -2633
rect 92 -2677 132 -2674
rect -386 -2689 -346 -2686
rect -386 -2723 -383 -2689
rect -349 -2723 -346 -2689
rect 92 -2711 95 -2677
rect 129 -2711 132 -2677
rect 2140 -2690 2240 -2667
rect 92 -2714 132 -2711
rect -386 -2726 -346 -2723
rect 2720 -2758 2830 -2750
rect 1870 -2773 2220 -2760
rect -248 -2826 106 -2778
rect 1870 -2807 2173 -2773
rect 2207 -2807 2220 -2773
rect 1870 -2810 2220 -2807
rect 1520 -2813 1560 -2810
rect 1520 -2847 1523 -2813
rect 1557 -2847 1560 -2813
rect 1880 -2830 2220 -2810
rect 2592 -2834 2830 -2758
rect 2720 -2840 2830 -2834
rect 1520 -2850 1560 -2847
rect -130 -2943 -50 -2910
rect -130 -2977 -107 -2943
rect -73 -2977 -50 -2943
rect -130 -3010 -50 -2977
rect 3070 -3080 3140 -1680
rect 2670 -3150 3140 -3080
<< viali >>
rect -187 -627 -153 -593
rect 2502 -662 2536 -628
rect 363 -787 397 -753
rect 2103 -817 2137 -783
rect -797 -947 -763 -913
rect -787 -1637 -753 -1603
rect 1703 -1787 1737 -1753
rect -635 -1851 -601 -1817
rect 2067 -1807 2101 -1773
rect -534 -1854 -500 -1820
rect 1024 -1952 1058 -1918
rect 1138 -1950 1172 -1916
rect -787 -1987 -753 -1953
rect 453 -2067 487 -2033
rect 1693 -2097 1727 -2063
rect 2173 -2667 2207 -2633
rect -383 -2723 -349 -2689
rect 95 -2711 129 -2677
rect 2173 -2807 2207 -2773
rect 1523 -2847 1557 -2813
rect 2424 -2942 2458 -2908
rect -107 -2977 -73 -2943
<< metal1 >>
rect -690 -530 -680 -440
rect -340 -540 0 -440
rect 1910 -540 2280 -440
rect -210 -593 -130 -540
rect -210 -627 -187 -593
rect -153 -627 -130 -593
rect -210 -660 -130 -627
rect 2490 -628 2950 -610
rect 2490 -662 2502 -628
rect 2536 -662 2950 -628
rect 2490 -680 2950 -662
rect -210 -753 420 -730
rect -210 -787 363 -753
rect 397 -787 420 -753
rect -210 -810 420 -787
rect 2080 -783 2150 -760
rect -820 -913 -740 -880
rect -820 -947 -797 -913
rect -763 -947 -740 -913
rect -820 -980 -740 -947
rect -820 -1080 -680 -980
rect -810 -1580 -660 -1480
rect -810 -1603 -730 -1580
rect -810 -1637 -787 -1603
rect -753 -1637 -730 -1603
rect -810 -1670 -730 -1637
rect -470 -1800 -380 -1790
rect -830 -1817 -580 -1800
rect -830 -1851 -635 -1817
rect -601 -1851 -580 -1817
rect -830 -1870 -580 -1851
rect -550 -1804 -380 -1800
rect -550 -1820 -446 -1804
rect -550 -1854 -534 -1820
rect -500 -1854 -446 -1820
rect -550 -1856 -446 -1854
rect -394 -1856 -380 -1804
rect -550 -1870 -380 -1856
rect -470 -1880 -380 -1870
rect -810 -1953 -730 -1920
rect -810 -1987 -787 -1953
rect -753 -1987 -730 -1953
rect -810 -2020 -730 -1987
rect -810 -2130 -670 -2020
rect -210 -2180 -140 -810
rect 2080 -817 2103 -783
rect 2137 -817 2150 -783
rect 730 -864 830 -840
rect 730 -916 754 -864
rect 806 -916 830 -864
rect 730 -930 830 -916
rect 440 -2033 510 -1070
rect 2080 -1330 2150 -817
rect 610 -1400 2150 -1330
rect 610 -1730 680 -1400
rect 1570 -1670 1850 -1570
rect 610 -1800 1190 -1730
rect 1000 -1918 1070 -1900
rect 1120 -1910 1190 -1800
rect 1680 -1753 1760 -1670
rect 1680 -1787 1703 -1753
rect 1737 -1787 1760 -1753
rect 1680 -1820 1760 -1787
rect 2050 -1773 2110 -1750
rect 2050 -1807 2067 -1773
rect 2101 -1807 2110 -1773
rect 2050 -1890 2110 -1807
rect 1000 -1952 1024 -1918
rect 1058 -1952 1070 -1918
rect 1000 -1970 1070 -1952
rect 1100 -1916 1210 -1910
rect 1100 -1950 1138 -1916
rect 1172 -1950 1210 -1916
rect 1100 -1960 1210 -1950
rect 2050 -1960 2280 -1890
rect 2050 -1962 2110 -1960
rect 440 -2067 453 -2033
rect 487 -2067 510 -2033
rect 440 -2090 510 -2067
rect 610 -2040 1070 -1970
rect -740 -2240 -140 -2180
rect -740 -2670 -670 -2240
rect 610 -2380 680 -2040
rect 1660 -2063 1760 -2040
rect 1660 -2097 1693 -2063
rect 1727 -2097 1760 -2063
rect 1660 -2120 1760 -2097
rect 1570 -2220 1850 -2120
rect 2880 -2340 2950 -680
rect -140 -2450 680 -2380
rect 2010 -2410 2950 -2340
rect -140 -2660 -70 -2450
rect -740 -2689 -330 -2670
rect -740 -2723 -383 -2689
rect -349 -2723 -330 -2689
rect -740 -2740 -330 -2723
rect -140 -2677 150 -2660
rect -140 -2711 95 -2677
rect 129 -2711 150 -2677
rect -140 -2740 150 -2711
rect 1110 -2674 1210 -2650
rect 1110 -2726 1134 -2674
rect 1186 -2726 1210 -2674
rect 1110 -2750 1210 -2726
rect 1490 -2813 1570 -2780
rect 1490 -2847 1523 -2813
rect 1557 -2820 1570 -2813
rect 2010 -2820 2080 -2410
rect 2140 -2633 2240 -2610
rect 2140 -2667 2173 -2633
rect 2207 -2667 2240 -2633
rect 2140 -2690 2240 -2667
rect 1557 -2847 2080 -2820
rect 2150 -2773 2480 -2760
rect 2150 -2807 2173 -2773
rect 2207 -2807 2480 -2773
rect 2150 -2830 2480 -2807
rect 1490 -2880 2080 -2847
rect 1490 -2890 1730 -2880
rect 1850 -2890 2080 -2880
rect 2410 -2908 2480 -2830
rect -130 -2943 -50 -2910
rect -130 -2977 -107 -2943
rect -73 -2977 -50 -2943
rect -130 -3060 -50 -2977
rect 2410 -2942 2424 -2908
rect 2458 -2942 2480 -2908
rect 2410 -2990 2480 -2942
rect -230 -3150 10 -3060
rect 1920 -3150 2320 -3060
<< via1 >>
rect -446 -1856 -394 -1804
rect 754 -916 806 -864
rect 1134 -2726 1186 -2674
<< metal2 >>
rect 730 -864 830 -840
rect 730 -916 754 -864
rect 806 -916 830 -864
rect 730 -950 830 -916
rect 730 -1180 800 -950
rect 100 -1250 800 -1180
rect -470 -1800 -380 -1790
rect 100 -1800 170 -1250
rect -470 -1804 170 -1800
rect -470 -1856 -446 -1804
rect -394 -1856 170 -1804
rect -470 -1870 170 -1856
rect -470 -1880 -380 -1870
rect 100 -2260 170 -1870
rect 100 -2330 1180 -2260
rect 1110 -2650 1180 -2330
rect 1110 -2674 1210 -2650
rect 1110 -2726 1134 -2674
rect 1186 -2726 1210 -2674
rect 1110 -2750 1210 -2726
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1729593089
transform -1 0 2680 0 -1 -2562
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1729593089
transform 1 0 1846 0 1 -2168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1729593089
transform 1 0 2280 0 1 -1032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_4
timestamp 1729593089
transform 1 0 -702 0 1 -1032
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_0
timestamp 1729593089
transform 1 0 -14 0 1 -1032
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_1
timestamp 1729593089
transform -1 0 1926 0 -1 -2562
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1729593089
transform 1 0 -672 0 1 -2074
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1729593089
transform -1 0 -224 0 -1 -2562
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1729593089
transform 1 0 930 0 1 -2168
box -38 -48 682 592
<< labels >>
rlabel metal1 s 2770 -610 2770 -610 4 Q1_buf
rlabel locali s 2040 -840 2040 -840 4 Q1
rlabel locali s 1620 -1940 1620 -1940 4 Dout
rlabel metal1 s 850 -1970 850 -1970 4 Q2
rlabel metal1 s -210 -1140 -210 -1140 4 Q2N
rlabel metal2 s -330 -1800 -330 -1800 4 SetBi
rlabel locali s -280 -810 -280 -810 4 UP_buf
rlabel metal1 s 2260 -2760 2260 -2760 4 DWN_buf
rlabel locali s -770 -760 -770 -760 4 UP
rlabel metal1 s -780 -1800 -780 -1800 4 SetB
rlabel locali s 2780 -2750 2780 -2750 4 DOWN
rlabel metal1 s 2270 -1890 2270 -1890 4 Dout_buf
rlabel locali s -320 -2020 -320 -2020 4 GND
rlabel locali s 2790 -470 2790 -470 4 VCCD
<< end >>
