magic
tech sky130A
timestamp 1725445935
<< error_p >>
rect -65 -40 425 540
rect -40 -510 0 -110
rect 365 -510 405 -110
<< nwell >>
rect -65 -40 425 540
<< pwell >>
rect -60 -550 425 -70
<< nmos >>
rect 0 -510 365 -110
<< pmos >>
rect 0 0 365 500
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -320 0 -300
rect -40 -340 -30 -320
rect -10 -340 0 -320
rect -40 -360 0 -340
rect -40 -380 -30 -360
rect -10 -380 0 -360
rect -40 -400 0 -380
rect -40 -420 -30 -400
rect -10 -420 0 -400
rect -40 -440 0 -420
rect -40 -460 -30 -440
rect -10 -460 0 -440
rect -40 -480 0 -460
rect -40 -500 -30 -480
rect -10 -500 0 -480
rect -40 -510 0 -500
rect 365 -120 405 -110
rect 365 -140 375 -120
rect 395 -140 405 -120
rect 365 -160 405 -140
rect 365 -180 375 -160
rect 395 -180 405 -160
rect 365 -200 405 -180
rect 365 -220 375 -200
rect 395 -220 405 -200
rect 365 -240 405 -220
rect 365 -260 375 -240
rect 395 -260 405 -240
rect 365 -280 405 -260
rect 365 -300 375 -280
rect 395 -300 405 -280
rect 365 -320 405 -300
rect 365 -340 375 -320
rect 395 -340 405 -320
rect 365 -360 405 -340
rect 365 -380 375 -360
rect 395 -380 405 -360
rect 365 -400 405 -380
rect 365 -420 375 -400
rect 395 -420 405 -400
rect 365 -440 405 -420
rect 365 -460 375 -440
rect 395 -460 405 -440
rect 365 -480 405 -460
rect 365 -500 375 -480
rect 395 -500 405 -480
rect 365 -510 405 -500
<< pdiff >>
rect -40 490 0 500
rect -40 470 -30 490
rect -10 470 0 490
rect -40 450 0 470
rect -40 430 -30 450
rect -10 430 0 450
rect -40 410 0 430
rect -40 390 -30 410
rect -10 390 0 410
rect -40 370 0 390
rect -40 350 -30 370
rect -10 350 0 370
rect -40 330 0 350
rect -40 310 -30 330
rect -10 310 0 330
rect -40 290 0 310
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 365 490 405 500
rect 365 470 375 490
rect 395 470 405 490
rect 365 450 405 470
rect 365 430 375 450
rect 395 430 405 450
rect 365 410 405 430
rect 365 390 375 410
rect 395 390 405 410
rect 365 370 405 390
rect 365 350 375 370
rect 395 350 405 370
rect 365 330 405 350
rect 365 310 375 330
rect 395 310 405 330
rect 365 290 405 310
rect 365 270 375 290
rect 395 270 405 290
rect 365 250 405 270
rect 365 230 375 250
rect 395 230 405 250
rect 365 210 405 230
rect 365 190 375 210
rect 395 190 405 210
rect 365 170 405 190
rect 365 150 375 170
rect 395 150 405 170
rect 365 130 405 150
rect 365 110 375 130
rect 395 110 405 130
rect 365 90 405 110
rect 365 70 375 90
rect 395 70 405 90
rect 365 50 405 70
rect 365 30 375 50
rect 395 30 405 50
rect 365 0 405 30
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect -30 -340 -10 -320
rect -30 -380 -10 -360
rect -30 -420 -10 -400
rect -30 -460 -10 -440
rect -30 -500 -10 -480
rect 375 -140 395 -120
rect 375 -180 395 -160
rect 375 -220 395 -200
rect 375 -260 395 -240
rect 375 -300 395 -280
rect 375 -340 395 -320
rect 375 -380 395 -360
rect 375 -420 395 -400
rect 375 -460 395 -440
rect 375 -500 395 -480
<< pdiffc >>
rect -30 470 -10 490
rect -30 430 -10 450
rect -30 390 -10 410
rect -30 350 -10 370
rect -30 310 -10 330
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 375 470 395 490
rect 375 430 395 450
rect 375 390 395 410
rect 375 350 395 370
rect 375 310 395 330
rect 375 270 395 290
rect 375 230 395 250
rect 375 190 395 210
rect 375 150 395 170
rect 375 110 395 130
rect 375 70 395 90
rect 375 30 395 50
<< poly >>
rect 0 500 365 540
rect 0 -110 365 0
rect 0 -550 365 -510
<< locali >>
rect -40 490 0 500
rect -40 470 -30 490
rect -10 470 0 490
rect -40 450 0 470
rect -40 430 -30 450
rect -10 430 0 450
rect -40 410 0 430
rect -40 390 -30 410
rect -10 390 0 410
rect -40 370 0 390
rect -40 350 -30 370
rect -10 350 0 370
rect -40 330 0 350
rect -40 310 -30 330
rect -10 310 0 330
rect -40 290 0 310
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 365 490 405 500
rect 365 470 375 490
rect 395 470 405 490
rect 365 450 405 470
rect 365 430 375 450
rect 395 430 405 450
rect 365 410 405 430
rect 365 390 375 410
rect 395 390 405 410
rect 365 370 405 390
rect 365 350 375 370
rect 395 350 405 370
rect 365 330 405 350
rect 365 310 375 330
rect 395 310 405 330
rect 365 290 405 310
rect 365 270 375 290
rect 395 270 405 290
rect 365 250 405 270
rect 365 230 375 250
rect 395 230 405 250
rect 365 210 405 230
rect 365 190 375 210
rect 395 190 405 210
rect 365 170 405 190
rect 365 150 375 170
rect 395 150 405 170
rect 365 130 405 150
rect 365 110 375 130
rect 395 110 405 130
rect 365 90 405 110
rect 365 70 375 90
rect 395 70 405 90
rect 365 50 405 70
rect 365 30 375 50
rect 395 30 405 50
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -320 0 -300
rect -40 -340 -30 -320
rect -10 -340 0 -320
rect -40 -360 0 -340
rect -40 -380 -30 -360
rect -10 -380 0 -360
rect -40 -400 0 -380
rect -40 -420 -30 -400
rect -10 -420 0 -400
rect -40 -440 0 -420
rect -40 -460 -30 -440
rect -10 -460 0 -440
rect -40 -480 0 -460
rect -40 -500 -30 -480
rect -10 -500 0 -480
rect -40 -510 0 -500
rect 365 -120 405 30
rect 365 -140 375 -120
rect 395 -140 405 -120
rect 365 -160 405 -140
rect 365 -180 375 -160
rect 395 -180 405 -160
rect 365 -200 405 -180
rect 365 -220 375 -200
rect 395 -220 405 -200
rect 365 -240 405 -220
rect 365 -260 375 -240
rect 395 -260 405 -240
rect 365 -280 405 -260
rect 365 -300 375 -280
rect 395 -300 405 -280
rect 365 -320 405 -300
rect 365 -340 375 -320
rect 395 -340 405 -320
rect 365 -360 405 -340
rect 365 -380 375 -360
rect 395 -380 405 -360
rect 365 -400 405 -380
rect 365 -420 375 -400
rect 395 -420 405 -400
rect 365 -440 405 -420
rect 365 -460 375 -440
rect 395 -460 405 -440
rect 365 -480 405 -460
rect 365 -500 375 -480
rect 395 -500 405 -480
rect 365 -510 405 -500
<< labels >>
rlabel poly 0 -55 0 -55 7 A
port 1 w
rlabel locali -20 500 -20 500 1 VPWR
port 2 n
rlabel locali -20 -510 -20 -510 5 VGND
port 3 s
rlabel locali 405 -55 405 -55 3 Y
port 4 e
<< end >>
