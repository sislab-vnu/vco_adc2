magic
tech sky130A
timestamp 1723626483
<< error_p >>
rect -90 -20 190 350
rect -70 -280 0 -80
rect 100 -280 170 -80
<< nwell >>
rect -90 -20 190 350
<< pwell >>
rect -90 -310 190 -60
<< nmos >>
rect 0 -280 100 -80
<< pmos >>
rect 0 0 100 300
<< ndiff >>
rect -70 -100 0 -80
rect -70 -130 -50 -100
rect -20 -130 0 -100
rect -70 -160 0 -130
rect -70 -190 -50 -160
rect -20 -190 0 -160
rect -70 -220 0 -190
rect -70 -250 -50 -220
rect -20 -250 0 -220
rect -70 -280 0 -250
rect 100 -100 170 -80
rect 100 -130 120 -100
rect 150 -130 170 -100
rect 100 -160 170 -130
rect 100 -190 120 -160
rect 150 -190 170 -160
rect 100 -220 170 -190
rect 100 -250 120 -220
rect 150 -250 170 -220
rect 100 -280 170 -250
<< pdiff >>
rect -70 280 0 300
rect -70 250 -50 280
rect -20 250 0 280
rect -70 220 0 250
rect -70 190 -50 220
rect -20 190 0 220
rect -70 160 0 190
rect -70 130 -50 160
rect -20 130 0 160
rect -70 100 0 130
rect -70 70 -50 100
rect -20 70 0 100
rect -70 50 0 70
rect -70 20 -50 50
rect -20 20 0 50
rect -70 0 0 20
rect 100 280 170 300
rect 100 250 120 280
rect 150 250 170 280
rect 100 220 170 250
rect 100 190 120 220
rect 150 190 170 220
rect 100 160 170 190
rect 100 130 120 160
rect 150 130 170 160
rect 100 100 170 130
rect 100 70 120 100
rect 150 70 170 100
rect 100 50 170 70
rect 100 20 120 50
rect 150 20 170 50
rect 100 0 170 20
<< ndiffc >>
rect -50 -130 -20 -100
rect -50 -190 -20 -160
rect -50 -250 -20 -220
rect 120 -130 150 -100
rect 120 -190 150 -160
rect 120 -250 150 -220
<< pdiffc >>
rect -50 250 -20 280
rect -50 190 -20 220
rect -50 130 -20 160
rect -50 70 -20 100
rect -50 20 -20 50
rect 120 250 150 280
rect 120 190 150 220
rect 120 130 150 160
rect 120 70 150 100
rect 120 20 150 50
<< poly >>
rect 0 300 100 330
rect 0 -80 100 0
rect 0 -310 100 -280
<< locali >>
rect -70 280 0 300
rect -70 250 -50 280
rect -20 250 0 280
rect -70 220 0 250
rect -70 190 -50 220
rect -20 190 0 220
rect -70 160 0 190
rect -70 130 -50 160
rect -20 130 0 160
rect -70 100 0 130
rect -70 70 -50 100
rect -20 70 0 100
rect -70 50 0 70
rect -70 20 -50 50
rect -20 20 0 50
rect -70 0 0 20
rect 100 280 170 300
rect 100 250 120 280
rect 150 250 170 280
rect 100 220 170 250
rect 100 190 120 220
rect 150 190 170 220
rect 100 160 170 190
rect 100 130 120 160
rect 150 130 170 160
rect 100 100 170 130
rect 100 70 120 100
rect 150 70 170 100
rect 100 50 170 70
rect 100 20 120 50
rect 150 20 170 50
rect 100 0 170 20
rect -70 -100 0 -80
rect -70 -130 -50 -100
rect -20 -130 0 -100
rect -70 -160 0 -130
rect -70 -190 -50 -160
rect -20 -190 0 -160
rect -70 -220 0 -190
rect -70 -250 -50 -220
rect -20 -250 0 -220
rect -70 -280 0 -250
rect 100 -100 170 -80
rect 100 -130 120 -100
rect 150 -130 170 -100
rect 100 -160 170 -130
rect 100 -190 120 -160
rect 150 -190 170 -160
rect 100 -220 170 -190
rect 100 -250 120 -220
rect 150 -250 170 -220
rect 100 -280 170 -250
<< end >>
