* NGSPICE file created from cc_inv.ext - technology: sky130A

.subckt aux_inv A Y VGND VDDA GND
X0 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt main_inv A Y VGND GND VDDA
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt cc_inv inp inn outp outn VGND VDDA GND
Xaux_inv_0 outp outn VGND VDDA GND aux_inv
Xaux_inv_1 outn outp VGND VDDA GND aux_inv
Xmain_inv_0 inp outp VGND GND VDDA main_inv
Xmain_inv_1 inn outn VGND GND VDDA main_inv
.ends


