magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -410 310 20 640
rect 520 300 940 630
rect -610 -530 -440 -210
rect 180 -540 650 -210
rect 2640 -260 2940 -210
rect 2630 -270 2940 -260
rect 2640 -540 2940 -270
<< pwell >>
rect -376 74 -244 226
rect -576 -806 -444 -654
rect 2634 -746 2786 -614
<< psubdiff >>
rect -350 167 -270 200
rect -350 133 -327 167
rect -293 133 -270 167
rect -350 100 -270 133
rect 2660 -663 2760 -640
rect -550 -713 -470 -680
rect -550 -747 -527 -713
rect -493 -747 -470 -713
rect 2660 -697 2693 -663
rect 2727 -697 2760 -663
rect 2660 -720 2760 -697
rect -550 -780 -470 -747
<< nsubdiff >>
rect -350 497 -270 530
rect -350 463 -327 497
rect -293 463 -270 497
rect -350 430 -270 463
rect -550 -353 -470 -320
rect -550 -387 -527 -353
rect -493 -387 -470 -353
rect -550 -420 -470 -387
rect 2680 -433 2780 -410
rect 2680 -467 2713 -433
rect 2747 -467 2780 -433
rect 2680 -490 2780 -467
<< psubdiffcont >>
rect -327 133 -293 167
rect -527 -747 -493 -713
rect 2693 -697 2727 -663
<< nsubdiffcont >>
rect -327 463 -293 497
rect -527 -387 -493 -353
rect 2713 -467 2747 -433
<< locali >>
rect 2420 570 2690 640
rect -350 497 -270 530
rect -350 463 -327 497
rect -293 463 -270 497
rect -350 430 -270 463
rect 70 307 110 310
rect 70 273 73 307
rect 107 273 110 307
rect 470 290 980 370
rect 70 270 110 273
rect 1240 247 1280 250
rect 1240 213 1243 247
rect 1277 213 1280 247
rect 1240 210 1280 213
rect -880 167 -270 200
rect -880 133 -847 167
rect -813 133 -327 167
rect -293 133 -270 167
rect -880 100 -270 133
rect 680 167 790 200
rect 680 133 723 167
rect 757 133 790 167
rect 2350 187 2390 190
rect 2350 153 2353 187
rect 2387 153 2390 187
rect 2350 150 2390 153
rect 680 110 790 133
rect 715 -65 765 110
rect 560 -115 765 -65
rect 150 -223 480 -200
rect 150 -257 413 -223
rect 447 -257 480 -223
rect 150 -290 480 -257
rect -550 -353 -470 -320
rect -550 -387 -527 -353
rect -493 -387 -470 -353
rect 560 -370 610 -115
rect 2610 -123 2690 570
rect 2610 -157 2633 -123
rect 2667 -157 2690 -123
rect 2610 -180 2690 -157
rect -550 -420 -470 -387
rect 150 -420 610 -370
rect 2070 -353 2110 -350
rect 2070 -387 2073 -353
rect 2107 -387 2110 -353
rect 2070 -390 2110 -387
rect 150 -530 205 -420
rect 2070 -433 2110 -430
rect 2070 -467 2073 -433
rect 2107 -467 2110 -433
rect 2070 -470 2110 -467
rect 2680 -433 2780 -410
rect 2680 -467 2713 -433
rect 2747 -467 2780 -433
rect 2680 -490 2780 -467
rect -700 -570 -370 -530
rect -700 -1000 -640 -570
rect 0 -580 205 -530
rect 2490 -530 2500 -520
rect 710 -543 750 -540
rect 710 -577 713 -543
rect 747 -577 750 -543
rect 2490 -570 2900 -530
rect 710 -580 750 -577
rect 960 -573 1000 -570
rect 960 -607 963 -573
rect 997 -607 1000 -573
rect 2490 -580 2500 -570
rect 2630 -600 2900 -570
rect 960 -610 1000 -607
rect 2070 -643 2110 -640
rect 2070 -677 2073 -643
rect 2107 -677 2110 -643
rect 2070 -680 2110 -677
rect 2660 -663 2760 -640
rect -550 -713 -470 -680
rect -550 -747 -527 -713
rect -493 -747 -470 -713
rect 2660 -697 2693 -663
rect 2727 -697 2760 -663
rect 2660 -720 2760 -697
rect -550 -780 -470 -747
rect 150 -840 680 -740
rect 2820 -1000 2900 -600
rect -700 -1080 2900 -1000
<< viali >>
rect -327 463 -293 497
rect 73 273 107 307
rect 1243 213 1277 247
rect -847 133 -813 167
rect -327 133 -293 167
rect 723 133 757 167
rect 2353 153 2387 187
rect 413 -257 447 -223
rect -527 -387 -493 -353
rect 2633 -157 2667 -123
rect 2073 -387 2107 -353
rect 2073 -467 2107 -433
rect 2713 -467 2747 -433
rect 713 -577 747 -543
rect 963 -607 997 -573
rect 2073 -677 2107 -643
rect -527 -747 -493 -713
rect 2693 -697 2727 -663
<< metal1 >>
rect 490 540 980 640
rect -720 497 -270 530
rect -720 463 -327 497
rect -293 463 -270 497
rect -720 430 -270 463
rect -880 167 -780 200
rect -880 133 -847 167
rect -813 133 -780 167
rect -880 -680 -780 133
rect -720 -320 -620 430
rect -500 307 140 330
rect -500 273 73 307
rect 107 273 140 307
rect -500 270 140 273
rect -500 -70 -440 270
rect 60 250 140 270
rect 1210 247 1310 290
rect 1210 220 1243 247
rect 680 213 1243 220
rect 1277 213 1310 247
rect -350 167 -270 200
rect -350 133 -327 167
rect -293 133 -270 167
rect -350 100 -270 133
rect 680 167 1310 213
rect 680 133 723 167
rect 757 150 1310 167
rect 2340 187 3330 230
rect 2340 153 2353 187
rect 2387 153 3330 187
rect 757 133 790 150
rect 680 110 790 133
rect 2340 130 3330 153
rect 490 0 960 70
rect 2430 0 3090 80
rect -500 -130 290 -70
rect -720 -353 -470 -320
rect -720 -387 -527 -353
rect -493 -387 -470 -353
rect -720 -420 -470 -387
rect 230 -540 290 -130
rect 2610 -123 2690 -100
rect 2610 -157 2633 -123
rect 2667 -157 2690 -123
rect 380 -223 690 -200
rect 380 -257 413 -223
rect 447 -257 690 -223
rect 380 -290 690 -257
rect 2610 -300 2690 -157
rect 2760 -330 2860 -130
rect 2050 -353 2860 -330
rect 2050 -387 2073 -353
rect 2107 -380 2860 -353
rect 2107 -387 2140 -380
rect 2050 -433 2140 -387
rect 2050 -467 2073 -433
rect 2107 -467 2140 -433
rect 690 -540 770 -470
rect 230 -543 770 -540
rect 230 -577 713 -543
rect 747 -577 770 -543
rect 230 -600 770 -577
rect 950 -573 1030 -530
rect 950 -607 963 -573
rect 997 -607 1030 -573
rect 950 -650 1030 -607
rect -880 -713 -470 -680
rect -880 -747 -527 -713
rect -493 -747 -470 -713
rect -880 -780 -470 -747
rect 480 -700 1030 -650
rect 2050 -540 2140 -467
rect 2680 -433 2780 -410
rect 2680 -467 2713 -433
rect 2747 -467 2780 -433
rect 2680 -490 2780 -467
rect 2050 -643 2150 -540
rect 2050 -677 2073 -643
rect 2107 -677 2150 -643
rect 2050 -690 2150 -677
rect 2660 -663 2760 -640
rect 2660 -697 2693 -663
rect 2727 -697 2760 -663
rect 480 -1150 580 -700
rect 2660 -720 2760 -697
rect 3000 -750 3090 0
rect 2610 -840 3090 -750
rect 3230 -1150 3330 130
rect 480 -1250 3330 -1150
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0
timestamp 1729593089
transform 1 0 -402 0 1 -792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_2  sky130_fd_sc_hd__dfxbp_2_0
timestamp 1729593089
transform 1 0 678 0 1 -792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1729593089
transform 1 0 958 0 1 48
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1729593089
transform 1 0 38 0 1 48
box -38 -48 498 592
<< labels >>
rlabel locali s 180 -580 180 -580 4 Q_N_buf
rlabel locali s -660 -530 -660 -530 4 Q_N
rlabel metal1 s 2580 230 2580 230 4 D
rlabel metal1 s -830 200 -830 200 4 VNB
rlabel metal1 s -510 530 -510 530 4 VPB
rlabel metal1 s 660 0 660 0 4 VGND
rlabel metal1 s 660 640 660 640 4 VPWR
rlabel locali s 680 290 680 290 4 clkinv
rlabel metal1 s 230 -70 230 -70 4 clk
rlabel metal1 s 2810 -130 2810 -130 4 clkDiv2
<< end >>
