magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -260 -80 600 680
<< pwell >>
rect -106 -504 586 -194
rect -246 -646 586 -504
rect -246 -656 -114 -646
<< nmos >>
rect 0 -620 200 -220
rect 280 -620 480 -220
<< pmos >>
rect 0 0 200 600
rect 280 0 480 600
<< ndiff >>
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -620 0 -597
rect 200 -243 280 -220
rect 200 -277 223 -243
rect 257 -277 280 -243
rect 200 -323 280 -277
rect 200 -357 223 -323
rect 257 -357 280 -323
rect 200 -403 280 -357
rect 200 -437 223 -403
rect 257 -437 280 -403
rect 200 -483 280 -437
rect 200 -517 223 -483
rect 257 -517 280 -483
rect 200 -563 280 -517
rect 200 -597 223 -563
rect 257 -597 280 -563
rect 200 -620 280 -597
rect 480 -243 560 -220
rect 480 -277 503 -243
rect 537 -277 560 -243
rect 480 -323 560 -277
rect 480 -357 503 -323
rect 537 -357 560 -323
rect 480 -403 560 -357
rect 480 -437 503 -403
rect 537 -437 560 -403
rect 480 -483 560 -437
rect 480 -517 503 -483
rect 537 -517 560 -483
rect 480 -563 560 -517
rect 480 -597 503 -563
rect 537 -597 560 -563
rect 480 -620 560 -597
<< pdiff >>
rect -80 577 0 600
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 200 577 280 600
rect 200 543 223 577
rect 257 543 280 577
rect 200 497 280 543
rect 200 463 223 497
rect 257 463 280 497
rect 200 417 280 463
rect 200 383 223 417
rect 257 383 280 417
rect 200 337 280 383
rect 200 303 223 337
rect 257 303 280 337
rect 200 257 280 303
rect 200 223 223 257
rect 257 223 280 257
rect 200 177 280 223
rect 200 143 223 177
rect 257 143 280 177
rect 200 97 280 143
rect 200 63 223 97
rect 257 63 280 97
rect 200 0 280 63
rect 480 577 560 600
rect 480 543 503 577
rect 537 543 560 577
rect 480 497 560 543
rect 480 463 503 497
rect 537 463 560 497
rect 480 417 560 463
rect 480 383 503 417
rect 537 383 560 417
rect 480 337 560 383
rect 480 303 503 337
rect 537 303 560 337
rect 480 257 560 303
rect 480 223 503 257
rect 537 223 560 257
rect 480 177 560 223
rect 480 143 503 177
rect 537 143 560 177
rect 480 97 560 143
rect 480 63 503 97
rect 537 63 560 97
rect 480 0 560 63
<< ndiffc >>
rect -57 -277 -23 -243
rect -57 -357 -23 -323
rect -57 -437 -23 -403
rect -57 -517 -23 -483
rect -57 -597 -23 -563
rect 223 -277 257 -243
rect 223 -357 257 -323
rect 223 -437 257 -403
rect 223 -517 257 -483
rect 223 -597 257 -563
rect 503 -277 537 -243
rect 503 -357 537 -323
rect 503 -437 537 -403
rect 503 -517 537 -483
rect 503 -597 537 -563
<< pdiffc >>
rect -57 543 -23 577
rect -57 463 -23 497
rect -57 383 -23 417
rect -57 303 -23 337
rect -57 223 -23 257
rect -57 143 -23 177
rect -57 63 -23 97
rect 223 543 257 577
rect 223 463 257 497
rect 223 383 257 417
rect 223 303 257 337
rect 223 223 257 257
rect 223 143 257 177
rect 223 63 257 97
rect 503 543 537 577
rect 503 463 537 497
rect 503 383 537 417
rect 503 303 537 337
rect 503 223 537 257
rect 503 143 537 177
rect 503 63 537 97
<< psubdiff >>
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
<< nsubdiff >>
rect -220 577 -140 610
rect -220 543 -197 577
rect -163 543 -140 577
rect -220 510 -140 543
<< psubdiffcont >>
rect -197 -597 -163 -563
<< nsubdiffcont >>
rect -197 543 -163 577
<< poly >>
rect 0 600 200 680
rect 280 600 480 680
rect 0 -80 200 0
rect 280 -80 480 0
rect 0 -93 480 -80
rect 0 -127 73 -93
rect 107 -127 363 -93
rect 397 -127 480 -93
rect 0 -140 480 -127
rect 0 -220 200 -140
rect 280 -220 480 -140
rect 0 -700 200 -620
rect 280 -700 480 -620
<< polycont >>
rect 73 -127 107 -93
rect 363 -127 397 -93
<< locali >>
rect -80 780 560 860
rect -220 577 -140 610
rect -220 543 -197 577
rect -163 543 -140 577
rect -220 510 -140 543
rect -80 577 0 780
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 200 577 280 600
rect 200 543 223 577
rect 257 543 280 577
rect 200 497 280 543
rect 200 463 223 497
rect 257 463 280 497
rect 200 417 280 463
rect 200 383 223 417
rect 257 383 280 417
rect 200 337 280 383
rect 200 303 223 337
rect 257 303 280 337
rect 200 257 280 303
rect 200 223 223 257
rect 257 223 280 257
rect 200 177 280 223
rect 200 143 223 177
rect 257 143 280 177
rect 200 97 280 143
rect 200 63 223 97
rect 257 63 280 97
rect 50 -93 140 -70
rect 50 -127 73 -93
rect 107 -127 140 -93
rect 50 -160 140 -127
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -800 0 -597
rect 200 -243 280 63
rect 480 577 560 780
rect 480 543 503 577
rect 537 543 560 577
rect 480 497 560 543
rect 480 463 503 497
rect 537 463 560 497
rect 480 417 560 463
rect 480 383 503 417
rect 537 383 560 417
rect 480 337 560 383
rect 480 303 503 337
rect 537 303 560 337
rect 480 257 560 303
rect 480 223 503 257
rect 537 223 560 257
rect 480 177 560 223
rect 480 143 503 177
rect 537 143 560 177
rect 480 97 560 143
rect 480 63 503 97
rect 537 63 560 97
rect 480 0 560 63
rect 330 -93 420 -70
rect 330 -127 363 -93
rect 397 -127 420 -93
rect 330 -160 420 -127
rect 200 -277 223 -243
rect 257 -277 280 -243
rect 200 -323 280 -277
rect 200 -357 223 -323
rect 257 -357 280 -323
rect 200 -403 280 -357
rect 200 -437 223 -403
rect 257 -437 280 -403
rect 200 -483 280 -437
rect 200 -517 223 -483
rect 257 -517 280 -483
rect 200 -563 280 -517
rect 200 -597 223 -563
rect 257 -597 280 -563
rect 200 -620 280 -597
rect 480 -243 560 -220
rect 480 -277 503 -243
rect 537 -277 560 -243
rect 480 -323 560 -277
rect 480 -357 503 -323
rect 537 -357 560 -323
rect 480 -403 560 -357
rect 480 -437 503 -403
rect 537 -437 560 -403
rect 480 -483 560 -437
rect 480 -517 503 -483
rect 537 -517 560 -483
rect 480 -563 560 -517
rect 480 -597 503 -563
rect 537 -597 560 -563
rect 480 -800 560 -597
rect -80 -880 560 -800
<< viali >>
rect -197 543 -163 577
rect 73 -127 107 -93
rect -197 -597 -163 -563
rect 363 -127 397 -93
<< metal1 >>
rect -220 577 -140 610
rect -220 543 -197 577
rect -163 543 -140 577
rect -220 510 -140 543
rect 50 -93 420 -70
rect 50 -127 73 -93
rect 107 -127 363 -93
rect 397 -127 420 -93
rect 50 -160 420 -127
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
<< labels >>
rlabel locali s 240 860 240 860 4 VPWR
rlabel metal1 s -180 610 -180 610 4 VCCA
rlabel locali s 240 600 240 600 4 Y
rlabel metal1 s -180 -530 -180 -530 4 GND
rlabel locali s 240 -800 240 -800 4 VGND
rlabel metal1 s 50 -110 50 -110 4 A
<< end >>
