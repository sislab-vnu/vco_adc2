magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -260 -80 320 680
<< pwell >>
rect -106 -504 306 -194
rect -246 -646 306 -504
rect -246 -656 -114 -646
<< nmos >>
rect 0 -620 200 -220
<< pmos >>
rect 0 0 200 600
<< ndiff >>
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -620 0 -597
rect 200 -243 280 -220
rect 200 -277 223 -243
rect 257 -277 280 -243
rect 200 -323 280 -277
rect 200 -357 223 -323
rect 257 -357 280 -323
rect 200 -403 280 -357
rect 200 -437 223 -403
rect 257 -437 280 -403
rect 200 -483 280 -437
rect 200 -517 223 -483
rect 257 -517 280 -483
rect 200 -563 280 -517
rect 200 -597 223 -563
rect 257 -597 280 -563
rect 200 -620 280 -597
<< pdiff >>
rect -80 577 0 600
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 200 577 280 600
rect 200 543 223 577
rect 257 543 280 577
rect 200 497 280 543
rect 200 463 223 497
rect 257 463 280 497
rect 200 417 280 463
rect 200 383 223 417
rect 257 383 280 417
rect 200 337 280 383
rect 200 303 223 337
rect 257 303 280 337
rect 200 257 280 303
rect 200 223 223 257
rect 257 223 280 257
rect 200 177 280 223
rect 200 143 223 177
rect 257 143 280 177
rect 200 97 280 143
rect 200 63 223 97
rect 257 63 280 97
rect 200 0 280 63
<< ndiffc >>
rect -57 -277 -23 -243
rect -57 -357 -23 -323
rect -57 -437 -23 -403
rect -57 -517 -23 -483
rect -57 -597 -23 -563
rect 223 -277 257 -243
rect 223 -357 257 -323
rect 223 -437 257 -403
rect 223 -517 257 -483
rect 223 -597 257 -563
<< pdiffc >>
rect -57 543 -23 577
rect -57 463 -23 497
rect -57 383 -23 417
rect -57 303 -23 337
rect -57 223 -23 257
rect -57 143 -23 177
rect -57 63 -23 97
rect 223 543 257 577
rect 223 463 257 497
rect 223 383 257 417
rect 223 303 257 337
rect 223 223 257 257
rect 223 143 257 177
rect 223 63 257 97
<< psubdiff >>
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
<< nsubdiff >>
rect -220 557 -140 590
rect -220 523 -197 557
rect -163 523 -140 557
rect -220 490 -140 523
<< psubdiffcont >>
rect -197 -597 -163 -563
<< nsubdiffcont >>
rect -197 523 -163 557
<< poly >>
rect 0 600 200 680
rect 0 -220 200 0
rect 0 -700 200 -620
<< locali >>
rect -220 557 -140 590
rect -220 523 -197 557
rect -163 523 -140 557
rect -220 490 -140 523
rect -80 577 0 600
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 200 577 280 600
rect 200 543 223 577
rect 257 543 280 577
rect 200 497 280 543
rect 200 463 223 497
rect 257 463 280 497
rect 200 417 280 463
rect 200 383 223 417
rect 257 383 280 417
rect 200 337 280 383
rect 200 303 223 337
rect 257 303 280 337
rect 200 257 280 303
rect 200 223 223 257
rect 257 223 280 257
rect 200 177 280 223
rect 200 143 223 177
rect 257 143 280 177
rect 200 97 280 143
rect 200 63 223 97
rect 257 63 280 97
rect -80 -243 0 -220
rect -80 -277 -57 -243
rect -23 -277 0 -243
rect -80 -323 0 -277
rect -80 -357 -57 -323
rect -23 -357 0 -323
rect -80 -403 0 -357
rect -80 -437 -57 -403
rect -23 -437 0 -403
rect -80 -483 0 -437
rect -80 -517 -57 -483
rect -23 -517 0 -483
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
rect -80 -563 0 -517
rect -80 -597 -57 -563
rect -23 -597 0 -563
rect -80 -620 0 -597
rect 200 -243 280 63
rect 200 -277 223 -243
rect 257 -277 280 -243
rect 200 -323 280 -277
rect 200 -357 223 -323
rect 257 -357 280 -323
rect 200 -403 280 -357
rect 200 -437 223 -403
rect 257 -437 280 -403
rect 200 -483 280 -437
rect 200 -517 223 -483
rect 257 -517 280 -483
rect 200 -563 280 -517
rect 200 -597 223 -563
rect 257 -597 280 -563
rect 200 -620 280 -597
<< viali >>
rect -197 523 -163 557
rect -197 -597 -163 -563
<< metal1 >>
rect -220 557 -140 590
rect -220 523 -197 557
rect -163 523 -140 557
rect -220 490 -140 523
rect -220 -563 -140 -530
rect -220 -597 -197 -563
rect -163 -597 -140 -563
rect -220 -630 -140 -597
<< labels >>
rlabel locali s -40 600 -40 600 4 VPWR
rlabel metal1 s -180 590 -180 590 4 VCCA
rlabel poly s 0 -110 0 -110 4 A
rlabel locali s 280 -110 280 -110 4 Y
rlabel metal1 s -180 -530 -180 -530 4 GND
rlabel locali s -40 -620 -40 -620 4 VGND
<< end >>
