* NGSPICE file created from aux_inv_vco.ext - technology: sky130A

.subckt nmos_vco_aux D G S VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt pmos_vco_aux D G S VPWR
X0 D G S VPWR sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
.ends

.subckt aux_inv_vco D G S_P S_N VPWR
Xnmos_vco_aux_0 D G S_N VSUBS nmos_vco_aux
Xpmos_vco_aux_0 D G S_P VPWR pmos_vco_aux
.ends

