** sch_path: /home/toind/work/vco_adc2/xschem/lib/vco_main_inv.sch
.subckt vco_main_inv VPWR VGND A Y VCCA GND
*.PININFO VPWR:B VGND:B A:I Y:O VCCA:B GND:B
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=3.65 W=8 nf=2 m=1
XM4 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 L=3.65 W=10 nf=2 m=1
.ends
.end
