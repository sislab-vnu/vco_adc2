magic
tech sky130A
timestamp 1726056110
<< nwell >>
rect 960 630 980 650
rect 960 590 980 610
<< pwell >>
rect 1250 260 1270 280
rect 1250 220 1270 240
<< ndiffc >>
rect 1250 260 1270 280
rect 1250 220 1270 240
<< pdiffc >>
rect 960 630 980 650
rect 960 590 980 610
<< polycont >>
rect 595 375 615 395
rect 885 375 905 395
<< locali >>
rect 335 830 1155 870
rect 520 740 560 830
rect 810 740 850 830
rect 585 395 625 405
rect 585 375 595 395
rect 615 375 625 395
rect 585 365 625 375
rect 700 395 915 405
rect 700 375 885 395
rect 905 375 915 395
rect 700 365 915 375
rect 520 40 560 130
rect 810 40 850 130
rect 300 0 1110 40
<< viali >>
rect 240 630 260 650
rect 960 630 980 650
rect 240 590 260 610
rect 960 590 980 610
rect 960 550 980 570
rect 670 470 690 490
rect 1250 470 1270 490
rect 595 375 615 395
rect 885 375 905 395
rect 1250 260 1270 280
rect 1250 220 1270 240
rect 1250 180 1270 200
<< metal1 >>
rect 20 950 1070 990
rect 20 745 60 950
rect 450 735 490 950
rect 740 735 780 950
rect 1030 745 1070 950
rect 230 650 270 660
rect 230 630 240 650
rect 260 640 270 650
rect 950 650 990 660
rect 950 640 960 650
rect 260 630 960 640
rect 980 630 990 650
rect 230 620 990 630
rect 0 580 195 620
rect 230 610 1440 620
rect 230 590 240 610
rect 260 600 960 610
rect 260 590 270 600
rect 230 580 270 590
rect 155 405 195 580
rect 585 395 625 600
rect 950 590 960 600
rect 980 590 1440 610
rect 950 580 1440 590
rect 950 570 990 580
rect 950 550 960 570
rect 980 550 990 570
rect 950 540 990 550
rect 660 490 1280 500
rect 660 470 670 490
rect 690 470 1250 490
rect 1270 470 1280 490
rect 660 460 1280 470
rect 585 375 595 395
rect 615 375 625 395
rect 585 365 625 375
rect 875 395 915 460
rect 875 375 885 395
rect 905 375 915 395
rect 875 365 915 375
rect 1165 250 1210 360
rect 0 210 1210 250
rect 1240 280 1280 290
rect 1240 260 1250 280
rect 1270 260 1280 280
rect 1240 250 1280 260
rect 1240 240 1440 250
rect 1240 220 1250 240
rect 1270 220 1440 240
rect 1240 210 1440 220
rect 1240 200 1280 210
rect 1240 180 1250 200
rect 1270 180 1280 200
rect 1240 170 1280 180
rect 20 -50 60 125
rect 450 -50 490 125
rect 740 -50 780 125
rect 1030 -50 1070 125
rect 20 -90 1070 -50
use dco_aux_inv  dco_aux_inv_0
timestamp 1726043895
transform 1 0 560 0 1 440
box -130 -350 160 340
use dco_aux_inv  dco_aux_inv_1
timestamp 1726043895
transform 1 0 850 0 1 440
box -130 -350 160 340
use dco_main_inv  dco_main_inv_0
timestamp 1726044335
transform 1 0 130 0 1 440
box -130 -440 300 430
use dco_main_inv  dco_main_inv_1
timestamp 1726044335
transform 1 0 1140 0 1 440
box -130 -440 300 430
<< labels >>
rlabel metal1 30 990 30 990 1 VCCA
port 1 n
rlabel metal1 0 600 0 600 7 inp
port 4 w
rlabel metal1 0 230 0 230 7 inn
port 5 w
rlabel metal1 65 -90 65 -90 5 GND
port 7 s
rlabel locali 645 870 645 870 1 VPWR
port 2 n
rlabel locali 655 0 655 0 5 VGND
port 8 s
rlabel metal1 1440 600 1440 600 3 outp
port 3 e
rlabel metal1 1440 230 1440 230 3 outn
port 6 e
<< end >>
