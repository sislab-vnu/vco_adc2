magic
tech sky130A
magscale 1 2
timestamp 1726657718
<< nwell >>
rect 380 220 420 260
rect 2220 220 2260 260
rect -690 -1760 -370 -1300
rect -680 -1810 -370 -1760
rect -690 -1860 -370 -1810
<< pwell >>
rect -930 -1780 -750 -1290
<< pdiffc >>
rect 380 220 420 260
rect 2220 220 2260 260
<< psubdiff >>
rect -890 -1640 -790 -1620
rect -890 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -890 -1700 -790 -1680
<< nsubdiff >>
rect -570 -1640 -470 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -470 -1640
rect -570 -1700 -470 -1680
<< psubdiffcont >>
rect -860 -1680 -820 -1640
<< nsubdiffcont >>
rect -540 -1680 -500 -1640
<< poly >>
rect 260 590 460 620
rect 260 550 360 590
rect 400 550 460 590
rect 2100 590 2300 620
rect 260 520 460 550
rect 2100 550 2200 590
rect 2240 550 2300 590
rect 2100 520 2300 550
<< polycont >>
rect 360 550 400 590
rect 1090 540 1130 580
rect 1210 540 1250 580
rect 1330 540 1370 580
rect 2200 550 2240 590
rect 2930 540 2970 580
rect 3050 540 3090 580
rect 3170 540 3210 580
<< locali >>
rect 160 940 850 1040
rect 180 450 260 830
rect 310 590 460 620
rect 310 550 360 590
rect 400 550 460 590
rect 310 520 460 550
rect 1040 580 1410 600
rect 1040 540 1090 580
rect 1130 540 1210 580
rect 1250 540 1330 580
rect 1370 540 1410 580
rect 1040 520 1410 540
rect 2150 590 2300 620
rect 2150 550 2200 590
rect 2240 550 2300 590
rect 2150 520 2300 550
rect 2880 580 3250 600
rect 2880 540 2930 580
rect 2970 540 3050 580
rect 3090 540 3170 580
rect 3210 540 3250 580
rect 2880 520 3250 540
rect 120 420 260 450
rect 120 350 180 420
rect 3300 -470 3380 110
rect 1020 -550 2110 -470
rect 2850 -550 3380 -470
rect -750 -980 -680 -770
rect -470 -1620 -360 -1290
rect -890 -1640 -790 -1620
rect -890 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -890 -1700 -790 -1680
rect -570 -1640 -360 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -440 -1640
rect -400 -1680 -360 -1640
rect -570 -1700 -360 -1680
rect -740 -1940 -690 -1930
rect -730 -2060 -690 -1940
rect -740 -2190 -690 -2060
rect -740 -2220 -620 -2190
rect -740 -2280 -710 -2220
rect -650 -2280 -620 -2220
rect -740 -2310 -620 -2280
rect 380 -2960 460 -2100
rect -1180 -3060 460 -2960
<< viali >>
rect 360 550 400 590
rect 1090 540 1130 580
rect 1210 540 1250 580
rect 1330 540 1370 580
rect 2200 550 2240 590
rect 2930 540 2970 580
rect 3050 540 3090 580
rect 3170 540 3210 580
rect 380 220 420 260
rect 2220 220 2260 260
rect 380 140 420 180
rect 2220 140 2260 180
rect -610 -1200 -570 -1160
rect -860 -1680 -820 -1640
rect -540 -1680 -500 -1640
rect -440 -1680 -400 -1640
rect -730 -1850 -690 -1810
rect -710 -2280 -650 -2220
<< metal1 >>
rect 1460 940 2840 1040
rect 260 590 460 620
rect 260 550 360 590
rect 400 550 460 590
rect 260 520 460 550
rect 1040 580 1410 600
rect 1040 540 1090 580
rect 1130 540 1210 580
rect 1250 540 1330 580
rect 1370 540 1410 580
rect 1040 520 1410 540
rect 360 260 440 280
rect 360 220 380 260
rect 420 220 440 260
rect 1460 240 1540 940
rect 2100 590 2300 620
rect 2100 550 2200 590
rect 2240 550 2300 590
rect 2100 520 2300 550
rect 2620 450 2700 940
rect 2760 440 2840 940
rect 2880 580 3250 600
rect 2880 540 2930 580
rect 2970 540 3050 580
rect 3090 540 3170 580
rect 3210 540 3250 580
rect 2880 520 3250 540
rect 360 180 440 220
rect 360 140 380 180
rect 420 140 440 180
rect 360 -60 440 140
rect 1880 -60 1960 400
rect 360 -140 1960 -60
rect 2200 260 2280 280
rect 2200 220 2220 260
rect 2260 220 2280 260
rect 2200 180 2280 220
rect 2200 140 2220 180
rect 2260 140 2280 180
rect 2200 -60 2280 140
rect 2200 -140 3530 -60
rect -230 -410 2830 -310
rect -1240 -620 -900 -520
rect -1000 -950 -900 -620
rect -999 -975 -904 -950
rect -760 -1160 -540 -1150
rect -760 -1200 -610 -1160
rect -570 -1200 -540 -1160
rect -760 -1210 -540 -1200
rect -1000 -1620 -900 -1310
rect -760 -1410 -680 -1210
rect -230 -1410 -130 -410
rect 380 -820 480 -410
rect -760 -1510 -130 -1410
rect 1770 -850 2250 -750
rect -1000 -1640 -790 -1620
rect -1000 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -1000 -1700 -790 -1680
rect -1000 -1780 -900 -1700
rect -760 -1810 -680 -1510
rect -570 -1640 -360 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -440 -1640
rect -400 -1680 -360 -1640
rect -570 -1700 -360 -1680
rect -470 -1780 -360 -1700
rect -760 -1850 -730 -1810
rect -690 -1850 -680 -1810
rect -760 -1870 -680 -1850
rect 1130 -2190 1250 -1510
rect 1770 -2190 1890 -850
rect 2730 -1480 2830 -410
rect 3450 -1320 3530 -140
rect 2730 -1560 3030 -1480
rect -740 -2220 1890 -2190
rect -740 -2280 -710 -2220
rect -650 -2280 1890 -2220
rect -740 -2310 1890 -2280
use obr  obr_0
timestamp 1726656757
transform 1 0 0 0 1 0
box 0 0 1580 1040
use obr  obr_1
timestamp 1726656757
transform 1 0 1840 0 1 0
box 0 0 1580 1040
use ol1  ol1_0
timestamp 1726656357
transform 1 0 20 0 1 -1810
box 0 -290 1580 1340
use ol1  ol1_1
timestamp 1726656357
transform 1 0 1990 0 1 -1810
box 0 -290 1580 1340
use sky130_fd_pr__res_xhigh_po_0p35_R469US  sky130_fd_pr__res_xhigh_po_0p35_R469US_0
timestamp 1726131431
transform -1 0 -1215 0 -1 -1788
box -35 -1272 35 1272
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 ~/eda/unic-cass/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -952 -1 0 -946
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 ~/eda/unic-cass/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -952 -1 0 -1776
box -38 -48 314 592
<< end >>
