magic
tech sky130A
magscale 1 2
timestamp 1730711120
<< locali >>
rect -2830 4030 3060 4050
rect -2830 3970 -2810 4030
rect -2750 3970 -2710 4030
rect -2650 3970 2740 4030
rect 2800 3970 2860 4030
rect 2920 3970 2980 4030
rect 3040 3970 3060 4030
rect -2830 3950 3060 3970
rect -2830 3930 -2730 3950
rect -2830 3870 -2810 3930
rect -2750 3870 -2730 3930
rect -2830 3850 -2730 3870
rect 2320 930 2420 3950
rect 2320 830 6030 930
rect 5930 -1180 6030 830
rect 5930 -1280 7040 -1180
rect 1130 -1560 6110 -1540
rect 1130 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 1130 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 6030 -1700 6110 -1680
rect 6940 -1690 7040 -1280
rect 6940 -1710 8290 -1690
rect 6940 -1770 8010 -1710
rect 8070 -1770 8110 -1710
rect 8170 -1770 8210 -1710
rect 8270 -1770 8290 -1710
rect 6940 -1790 8290 -1770
rect 1470 -2150 2740 -2130
rect 1470 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 1470 -2220 2740 -2210
rect 1530 -2230 2740 -2220
rect 1580 -2420 3950 -2400
rect 1580 -2480 3770 -2420
rect 3830 -2480 3870 -2420
rect 3930 -2480 3950 -2420
rect 1580 -2500 3950 -2480
rect 3850 -2520 3950 -2500
rect 3850 -2580 3870 -2520
rect 3930 -2580 3950 -2520
rect 3850 -2600 3950 -2580
rect 3850 -4790 3950 -4770
rect 3850 -4850 3870 -4790
rect 3930 -4850 3950 -4790
rect 3850 -4870 3950 -4850
rect 2080 -4890 3950 -4870
rect 2080 -4950 2100 -4890
rect 2160 -4950 2220 -4890
rect 2280 -4950 2340 -4890
rect 2400 -4950 3870 -4890
rect 3930 -4950 3950 -4890
rect 2080 -4970 3950 -4950
rect 3850 -4990 3950 -4970
rect 3850 -5050 3870 -4990
rect 3930 -5050 3950 -4990
rect 860 -5680 1060 -5050
rect 3850 -5070 3950 -5050
rect 860 -5720 880 -5680
rect 920 -5720 1000 -5680
rect 1040 -5720 1060 -5680
rect 860 -5810 1060 -5720
rect 860 -5850 880 -5810
rect 920 -5850 1000 -5810
rect 1040 -5850 1060 -5810
rect 860 -5870 1060 -5850
rect -2240 -6750 -1830 -6740
rect -2240 -6760 -1820 -6750
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -1820 -6760
rect -2240 -6820 -1820 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -2240 -6900 -2160 -6880
rect -2830 -7690 -2730 -7670
rect -2830 -7750 -2810 -7690
rect -2750 -7750 -2730 -7690
rect -2830 -7770 -2730 -7750
rect -2830 -7790 -1890 -7770
rect -2830 -7850 -2810 -7790
rect -2750 -7850 -2710 -7790
rect -2650 -7850 -2070 -7790
rect -2010 -7850 -1970 -7790
rect -1910 -7850 -1890 -7790
rect -2830 -7870 -1890 -7850
rect 1260 -7890 2370 -7870
rect 1260 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 1260 -7950 2370 -7930
rect 16280 -7900 17170 -7870
rect 16280 -7940 16310 -7900
rect 16350 -7940 16390 -7900
rect 16430 -7940 17170 -7900
rect 16280 -7970 17170 -7940
rect 16280 -7980 16380 -7970
rect 16280 -8020 16310 -7980
rect 16350 -8020 16380 -7980
rect 16280 -8050 16380 -8020
rect 3850 -8650 3950 -8630
rect 3850 -8710 3870 -8650
rect 3930 -8710 3950 -8650
rect 3850 -8730 3950 -8710
rect 1580 -8750 3950 -8730
rect 1580 -8810 3770 -8750
rect 3830 -8810 3870 -8750
rect 3930 -8810 3950 -8750
rect 1580 -8830 3950 -8810
rect -3060 -9140 -1540 -9080
rect -3060 -9220 -3020 -9140
rect -2940 -9220 -2860 -9140
rect -2780 -9220 -2700 -9140
rect -2620 -9220 -1540 -9140
rect -3060 -9280 -1540 -9220
rect 17070 -9960 17170 -7970
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect 17000 -10040 17170 -10020
rect 17000 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect 17000 -10100 17170 -10080
<< viali >>
rect -270 8010 -230 8050
rect -190 8010 -150 8050
rect -110 8010 -70 8050
rect -30 8010 10 8050
rect 50 8010 90 8050
rect 3040 8010 3080 8050
rect 3120 8010 3160 8050
rect 3200 8010 3240 8050
rect 3280 8010 3320 8050
rect 3360 8010 3400 8050
rect 11060 8010 11100 8050
rect 11140 8010 11180 8050
rect 11220 8010 11260 8050
rect 11300 8010 11340 8050
rect 11380 8010 11420 8050
rect 15890 8010 15930 8050
rect 15970 8010 16010 8050
rect 16050 8010 16090 8050
rect 16130 8010 16170 8050
rect 16210 8010 16250 8050
rect -2810 3970 -2750 4030
rect -2710 3970 -2650 4030
rect 2740 3970 2800 4030
rect 2860 3970 2920 4030
rect 2980 3970 3040 4030
rect -2810 3870 -2750 3930
rect -2000 -470 -1960 -430
rect -1920 -470 -1880 -430
rect 1150 -1600 1190 -1560
rect 1230 -1600 1270 -1560
rect 5970 -1600 6010 -1560
rect 6050 -1600 6090 -1560
rect 6050 -1680 6090 -1640
rect 8010 -1770 8070 -1710
rect 8110 -1770 8170 -1710
rect 8210 -1770 8270 -1710
rect 2420 -2210 2480 -2150
rect 2540 -2210 2600 -2150
rect 2660 -2210 2720 -2150
rect 3770 -2480 3830 -2420
rect 3870 -2480 3930 -2420
rect 3870 -2580 3930 -2520
rect 3870 -4850 3930 -4790
rect 2100 -4950 2160 -4890
rect 2220 -4950 2280 -4890
rect 2340 -4950 2400 -4890
rect 3870 -4950 3930 -4890
rect 3870 -5050 3930 -4990
rect 880 -5720 920 -5680
rect 1000 -5720 1040 -5680
rect 880 -5850 920 -5810
rect 1000 -5850 1040 -5810
rect -2220 -6800 -2180 -6760
rect -2140 -6800 -2100 -6760
rect -2220 -6880 -2180 -6840
rect -2810 -7750 -2750 -7690
rect -2810 -7850 -2750 -7790
rect -2710 -7850 -2650 -7790
rect -2070 -7850 -2010 -7790
rect -1970 -7850 -1910 -7790
rect 1280 -7930 1320 -7890
rect 1360 -7930 1400 -7890
rect 1440 -7930 1480 -7890
rect 2150 -7930 2190 -7890
rect 2230 -7930 2270 -7890
rect 2310 -7930 2350 -7890
rect 16310 -7940 16350 -7900
rect 16390 -7940 16430 -7900
rect 16310 -8020 16350 -7980
rect 3870 -8710 3930 -8650
rect 3770 -8810 3830 -8750
rect 3870 -8810 3930 -8750
rect -3020 -9220 -2940 -9140
rect -2860 -9220 -2780 -9140
rect -2700 -9220 -2620 -9140
rect 17100 -10000 17140 -9960
rect 17020 -10080 17060 -10040
rect 17100 -10080 17140 -10040
<< metal1 >>
rect -290 8060 110 8070
rect -290 8000 -280 8060
rect -220 8050 -160 8060
rect -100 8050 -40 8060
rect 20 8050 110 8060
rect -220 8010 -190 8050
rect -70 8010 -40 8050
rect 20 8010 50 8050
rect 90 8010 110 8050
rect -220 8000 -160 8010
rect -100 8000 -40 8010
rect 20 8000 110 8010
rect -290 7990 110 8000
rect 3020 8060 3420 8070
rect 3020 8000 3030 8060
rect 3090 8050 3190 8060
rect 3250 8050 3350 8060
rect 3090 8010 3120 8050
rect 3160 8010 3190 8050
rect 3250 8010 3280 8050
rect 3320 8010 3350 8050
rect 3090 8000 3190 8010
rect 3250 8000 3350 8010
rect 3410 8000 3420 8060
rect 3020 7990 3420 8000
rect 11040 8060 11440 8070
rect 11040 8000 11050 8060
rect 11110 8050 11210 8060
rect 11270 8050 11370 8060
rect 11110 8010 11140 8050
rect 11180 8010 11210 8050
rect 11270 8010 11300 8050
rect 11340 8010 11370 8050
rect 11110 8000 11210 8010
rect 11270 8000 11370 8010
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8060 16270 8070
rect 15870 8000 15880 8060
rect 15940 8050 16040 8060
rect 16100 8050 16200 8060
rect 15940 8010 15970 8050
rect 16010 8010 16040 8050
rect 16100 8010 16130 8050
rect 16170 8010 16200 8050
rect 15940 8000 16040 8010
rect 16100 8000 16200 8010
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 6900 4980 7140 5000
rect 6900 4920 6920 4980
rect 6980 4920 7040 4980
rect 7100 4920 7140 4980
rect 6900 4880 7140 4920
rect 6900 4820 6920 4880
rect 6980 4820 7040 4880
rect 7100 4820 7140 4880
rect 6900 4800 7140 4820
rect -2830 4030 -2630 4050
rect -2830 3970 -2810 4030
rect -2750 3970 -2710 4030
rect -2650 3970 -2630 4030
rect -2830 3930 -2630 3970
rect 2710 4030 3060 4050
rect 2710 3970 2740 4030
rect 2800 3970 2860 4030
rect 2920 3970 2980 4030
rect 3040 3970 3060 4030
rect 2710 3950 3060 3970
rect -2830 3870 -2810 3930
rect -2750 3870 -2630 3930
rect -2830 3770 -2630 3870
rect -2830 3670 -2790 3770
rect -2690 3670 -2630 3770
rect -2830 3570 -2630 3670
rect -2830 3470 -2790 3570
rect -2690 3470 -2630 3570
rect -2830 3370 -2630 3470
rect -2830 3270 -2790 3370
rect -2690 3270 -2630 3370
rect -2830 -1430 -2630 3270
rect -2020 -410 -1920 2100
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 -130 -1080 1010
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 -120 80 1000
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 -130 1290 1020
rect -2020 -430 -1860 -410
rect -2020 -470 -2000 -430
rect -1960 -470 -1920 -430
rect -1880 -470 -1860 -430
rect -2020 -490 -1860 -470
rect -2830 -1456 -2000 -1430
rect -2830 -1526 -1875 -1456
rect -2830 -1530 -2000 -1526
rect -2830 -7690 -2630 -1530
rect 970 -1560 1290 -1540
rect 970 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 1290 -1560
rect 970 -1620 1290 -1600
rect 5950 -1560 6110 -1540
rect 5950 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 5950 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 2400 -2150 2740 -2130
rect 2400 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 2400 -2230 2740 -2210
rect 2360 -3100 2760 -2230
rect 3750 -2420 3950 -2400
rect 3750 -2480 3770 -2420
rect 3830 -2480 3870 -2420
rect 3930 -2480 3950 -2420
rect 3750 -2500 3950 -2480
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3480 2760 -3280
rect 3850 -2520 3950 -2500
rect 3850 -2580 3870 -2520
rect 3930 -2580 3950 -2520
rect -2320 -4490 -1920 -3900
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4800 -1920 -4550
rect -1770 -4210 -1570 -4190
rect -1770 -4310 -1730 -4210
rect -1630 -4310 -1570 -4210
rect -1770 -4380 -1570 -4310
rect -1770 -4480 -1730 -4380
rect -1630 -4480 -1570 -4380
rect -1770 -4540 -1570 -4480
rect -1770 -4640 -1730 -4540
rect -1630 -4640 -1570 -4540
rect -1770 -4660 -1570 -4640
rect 3850 -4790 3950 -2580
rect 3850 -4850 3870 -4790
rect 3930 -4850 3950 -4790
rect 2080 -4890 2420 -4870
rect 2080 -4950 2100 -4890
rect 2160 -4950 2220 -4890
rect 2280 -4950 2340 -4890
rect 2400 -4950 2420 -4890
rect 2080 -4970 2420 -4950
rect 3850 -4890 3950 -4850
rect 3850 -4950 3870 -4890
rect 3930 -4950 3950 -4890
rect 6030 -4830 6110 -1680
rect 7990 -1710 8290 -1690
rect 7990 -1770 8010 -1710
rect 8070 -1770 8110 -1710
rect 8170 -1770 8210 -1710
rect 8270 -1770 8290 -1710
rect 7990 -1790 8290 -1770
rect 13160 -3580 13250 -3540
rect 13160 -3640 13170 -3580
rect 13230 -3640 13250 -3580
rect 13160 -3700 13250 -3640
rect 13160 -3760 13170 -3700
rect 13230 -3760 13250 -3700
rect 13160 -3890 13250 -3760
rect 6540 -4480 6740 -4460
rect 6540 -4540 6560 -4480
rect 6620 -4540 6660 -4480
rect 6720 -4500 6740 -4480
rect 6720 -4540 8190 -4500
rect 6540 -4580 8190 -4540
rect 6540 -4640 6560 -4580
rect 6620 -4640 6660 -4580
rect 6720 -4600 8190 -4580
rect 6720 -4640 6740 -4600
rect 6540 -4660 6740 -4640
rect 6030 -4910 6520 -4830
rect 3850 -4990 3950 -4950
rect -1790 -6070 -1710 -5020
rect 3850 -5050 3870 -4990
rect 3930 -5050 3950 -4990
rect -1480 -5500 -1080 -5340
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5580 -1080 -5560
rect -90 -5500 310 -5340
rect -90 -5560 -60 -5500
rect 0 -5560 60 -5500
rect 120 -5560 180 -5500
rect 240 -5560 310 -5500
rect -90 -5580 310 -5560
rect 860 -5680 1280 -5670
rect 860 -5720 880 -5680
rect 920 -5720 1000 -5680
rect 1040 -5690 1280 -5680
rect 1040 -5720 1080 -5690
rect 860 -5750 1080 -5720
rect 1140 -5750 1200 -5690
rect 1260 -5750 1280 -5690
rect 860 -5790 1280 -5750
rect 860 -5810 1080 -5790
rect 860 -5850 880 -5810
rect 920 -5850 1000 -5810
rect 1040 -5850 1080 -5810
rect 1140 -5850 1200 -5790
rect 1260 -5850 1280 -5790
rect 860 -5870 1280 -5850
rect -1790 -6150 2370 -6070
rect -2830 -7750 -2810 -7690
rect -2750 -7750 -2630 -7690
rect -2830 -7790 -2630 -7750
rect -2830 -7850 -2810 -7790
rect -2750 -7850 -2710 -7790
rect -2650 -7850 -2630 -7790
rect -2830 -7870 -2630 -7850
rect -2240 -6760 -2080 -6740
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -2080 -6760
rect -2240 -6820 -2080 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -3060 -9140 -2580 -9080
rect -3060 -9220 -3020 -9140
rect -2940 -9220 -2860 -9140
rect -2780 -9220 -2700 -9140
rect -2620 -9220 -2580 -9140
rect -3060 -9280 -2580 -9220
rect -3060 -9390 -2660 -9280
rect -3060 -9450 -3030 -9390
rect -2970 -9450 -2910 -9390
rect -2850 -9450 -2790 -9390
rect -2730 -9450 -2660 -9390
rect -3060 -9590 -2660 -9450
rect -2240 -10020 -2160 -6880
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7170 -1480 -7150
rect -2100 -7790 -1890 -7770
rect -2100 -7850 -2070 -7790
rect -2010 -7850 -1970 -7790
rect -1910 -7850 -1890 -7790
rect -2100 -7870 -1890 -7850
rect 2290 -7870 2370 -6150
rect 970 -7890 1500 -7870
rect 970 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 1500 -7890
rect 970 -7950 1500 -7930
rect 2130 -7890 2370 -7870
rect 2130 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 2130 -7950 2370 -7930
rect 3850 -8650 3950 -5050
rect 6440 -7010 6520 -4910
rect 9100 -4950 9300 -4930
rect 9100 -5010 9120 -4950
rect 9180 -5010 9220 -4950
rect 9280 -5010 9300 -4950
rect 9100 -5050 9300 -5010
rect 9100 -5110 9120 -5050
rect 9180 -5110 9220 -5050
rect 9280 -5110 9300 -5050
rect 9100 -5130 9300 -5110
rect 16280 -7900 16490 -7870
rect 16280 -7940 16310 -7900
rect 16350 -7940 16390 -7900
rect 16430 -7940 16490 -7900
rect 16280 -7970 16490 -7940
rect 16280 -7980 16380 -7970
rect 16280 -8020 16310 -7980
rect 16350 -8020 16380 -7980
rect 16280 -8050 16380 -8020
rect 12250 -8140 12650 -8120
rect 12250 -8200 12280 -8140
rect 12340 -8200 12400 -8140
rect 12460 -8200 12520 -8140
rect 12580 -8200 12650 -8140
rect 12250 -8220 12650 -8200
rect 3850 -8710 3870 -8650
rect 3930 -8710 3950 -8650
rect 3850 -8730 3950 -8710
rect 3750 -8750 3950 -8730
rect 3750 -8810 3770 -8750
rect 3830 -8810 3870 -8750
rect 3930 -8810 3950 -8750
rect 3750 -8830 3950 -8810
rect -1640 -9140 -1240 -9050
rect 580 -9160 980 -9060
rect 580 -9220 610 -9160
rect 670 -9220 730 -9160
rect 790 -9220 850 -9160
rect 910 -9220 980 -9160
rect 580 -9250 980 -9220
rect 17070 -9960 17170 -9940
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect -2240 -10040 17170 -10020
rect -2240 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect -2240 -10100 17170 -10080
<< via1 >>
rect -280 8050 -220 8060
rect -160 8050 -100 8060
rect -40 8050 20 8060
rect -280 8010 -270 8050
rect -270 8010 -230 8050
rect -230 8010 -220 8050
rect -160 8010 -150 8050
rect -150 8010 -110 8050
rect -110 8010 -100 8050
rect -40 8010 -30 8050
rect -30 8010 10 8050
rect 10 8010 20 8050
rect -280 8000 -220 8010
rect -160 8000 -100 8010
rect -40 8000 20 8010
rect 3030 8050 3090 8060
rect 3190 8050 3250 8060
rect 3350 8050 3410 8060
rect 3030 8010 3040 8050
rect 3040 8010 3080 8050
rect 3080 8010 3090 8050
rect 3190 8010 3200 8050
rect 3200 8010 3240 8050
rect 3240 8010 3250 8050
rect 3350 8010 3360 8050
rect 3360 8010 3400 8050
rect 3400 8010 3410 8050
rect 3030 8000 3090 8010
rect 3190 8000 3250 8010
rect 3350 8000 3410 8010
rect 11050 8050 11110 8060
rect 11210 8050 11270 8060
rect 11370 8050 11430 8060
rect 11050 8010 11060 8050
rect 11060 8010 11100 8050
rect 11100 8010 11110 8050
rect 11210 8010 11220 8050
rect 11220 8010 11260 8050
rect 11260 8010 11270 8050
rect 11370 8010 11380 8050
rect 11380 8010 11420 8050
rect 11420 8010 11430 8050
rect 11050 8000 11110 8010
rect 11210 8000 11270 8010
rect 11370 8000 11430 8010
rect 15880 8050 15940 8060
rect 16040 8050 16100 8060
rect 16200 8050 16260 8060
rect 15880 8010 15890 8050
rect 15890 8010 15930 8050
rect 15930 8010 15940 8050
rect 16040 8010 16050 8050
rect 16050 8010 16090 8050
rect 16090 8010 16100 8050
rect 16200 8010 16210 8050
rect 16210 8010 16250 8050
rect 16250 8010 16260 8050
rect 15880 8000 15940 8010
rect 16040 8000 16100 8010
rect 16200 8000 16260 8010
rect 6920 4920 6980 4980
rect 7040 4920 7100 4980
rect 6920 4820 6980 4880
rect 7040 4820 7100 4880
rect 14700 4500 14760 4560
rect 14700 4380 14760 4440
rect 14700 4260 14760 4320
rect -2790 3670 -2690 3770
rect -2790 3470 -2690 3570
rect -2790 3270 -2690 3370
rect -1430 1010 -1360 1080
rect -1200 1010 -1130 1080
rect -270 1000 -200 1070
rect -50 1000 20 1070
rect 930 1020 990 1080
rect 1180 1020 1240 1080
rect 2390 -3160 2450 -3100
rect 2510 -3160 2570 -3100
rect 2630 -3160 2690 -3100
rect 2390 -3280 2450 -3220
rect 2510 -3280 2570 -3220
rect 2630 -3280 2690 -3220
rect -2280 -4550 -2220 -4490
rect -2030 -4550 -1970 -4490
rect -1730 -4310 -1630 -4210
rect -1730 -4480 -1630 -4380
rect -1730 -4640 -1630 -4540
rect 18530 -2080 18590 -2020
rect 18530 -2200 18590 -2140
rect 18530 -2320 18590 -2260
rect 13170 -3640 13230 -3580
rect 13170 -3760 13230 -3700
rect 6560 -4540 6620 -4480
rect 6660 -4540 6720 -4480
rect 6560 -4640 6620 -4580
rect 6660 -4640 6720 -4580
rect -1450 -5560 -1390 -5500
rect -1330 -5560 -1270 -5500
rect -1210 -5560 -1150 -5500
rect -60 -5560 0 -5500
rect 60 -5560 120 -5500
rect 180 -5560 240 -5500
rect 1080 -5750 1140 -5690
rect 1200 -5750 1260 -5690
rect 1080 -5850 1140 -5790
rect 1200 -5850 1260 -5790
rect -3030 -9450 -2970 -9390
rect -2910 -9450 -2850 -9390
rect -2790 -9450 -2730 -9390
rect -1930 -7150 -1870 -7090
rect -1810 -7150 -1750 -7090
rect -1690 -7150 -1630 -7090
rect -1570 -7150 -1510 -7090
rect 9120 -5010 9180 -4950
rect 9220 -5010 9280 -4950
rect 9120 -5110 9180 -5050
rect 9220 -5110 9280 -5050
rect 18530 -7070 18590 -7010
rect 18530 -7190 18590 -7130
rect 18530 -7310 18590 -7250
rect 12280 -8200 12340 -8140
rect 12400 -8200 12460 -8140
rect 12520 -8200 12580 -8140
rect 610 -9220 670 -9160
rect 730 -9220 790 -9160
rect 850 -9220 910 -9160
rect 8030 -9640 8090 -9580
rect 8150 -9640 8210 -9580
rect 8270 -9640 8330 -9580
rect 16090 -9640 16150 -9580
rect 16210 -9640 16270 -9580
rect 16330 -9640 16390 -9580
<< metal2 >>
rect 17342 35320 17710 36938
rect 17342 34920 24990 35320
rect 17342 34914 17710 34920
rect -290 8180 110 8210
rect -290 8100 -250 8180
rect -170 8100 -10 8180
rect 70 8100 110 8180
rect -290 8060 110 8100
rect -290 8000 -280 8060
rect -220 8000 -160 8060
rect -100 8000 -40 8060
rect 20 8000 110 8060
rect -290 7990 110 8000
rect 3020 8190 3420 8210
rect 3020 8110 3060 8190
rect 3140 8110 3280 8190
rect 3360 8110 3420 8190
rect 3020 8060 3420 8110
rect 3020 8000 3030 8060
rect 3090 8000 3190 8060
rect 3250 8000 3350 8060
rect 3410 8000 3420 8060
rect 3020 7990 3420 8000
rect 11040 8190 11440 8220
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8060 11440 8110
rect 11040 8000 11050 8060
rect 11110 8000 11210 8060
rect 11270 8000 11370 8060
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8180 16270 8210
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8060 16270 8100
rect 15870 8000 15880 8060
rect 15940 8000 16040 8060
rect 16100 8000 16200 8060
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 24590 5000 24990 34920
rect 6900 4980 24990 5000
rect 6900 4920 6920 4980
rect 6980 4920 7040 4980
rect 7100 4920 24990 4980
rect 6900 4880 24990 4920
rect 6900 4820 6920 4880
rect 6980 4820 7040 4880
rect 7100 4820 24990 4880
rect 6900 4800 24990 4820
rect 14680 4570 14990 4630
rect 14680 4560 14830 4570
rect 14680 4500 14700 4560
rect 14760 4500 14830 4560
rect 14680 4470 14830 4500
rect 14930 4470 14990 4570
rect 14680 4440 14990 4470
rect 14680 4380 14700 4440
rect 14760 4380 14990 4440
rect 14680 4370 14990 4380
rect 14680 4320 14830 4370
rect 14680 4260 14700 4320
rect 14760 4270 14830 4320
rect 14930 4270 14990 4370
rect 14760 4260 14990 4270
rect 14680 4230 14990 4260
rect -7520 3770 -2630 3850
rect -7520 3670 -2790 3770
rect -2690 3670 -2630 3770
rect -7520 3570 -2630 3670
rect -7520 3470 -2790 3570
rect -2690 3470 -2630 3570
rect -7520 3450 -2630 3470
rect -7520 -17770 -7120 3450
rect -2830 3370 -2630 3450
rect -2830 3270 -2790 3370
rect -2690 3270 -2630 3370
rect -2830 3250 -2630 3270
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 960 -1080 1010
rect -1480 880 -1430 960
rect -1350 880 -1220 960
rect -1140 880 -1080 960
rect -1480 820 -1080 880
rect -1480 740 -1430 820
rect -1350 740 -1220 820
rect -1140 740 -1080 820
rect -1480 710 -1080 740
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 950 80 1000
rect -320 870 -270 950
rect -190 870 -50 950
rect 30 870 80 950
rect -320 810 80 870
rect -320 730 -270 810
rect -190 730 -50 810
rect 30 730 80 810
rect -320 710 80 730
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 980 1290 1020
rect 890 900 930 980
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 890 820 1290 900
rect 890 740 930 820
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 890 710 1290 740
rect 18510 -2000 18790 -1950
rect 18510 -2020 18650 -2000
rect 18510 -2080 18530 -2020
rect 18590 -2080 18650 -2020
rect 18730 -2080 18790 -2000
rect 18510 -2140 18790 -2080
rect 18510 -2200 18530 -2140
rect 18590 -2160 18790 -2140
rect 18590 -2200 18650 -2160
rect 18510 -2240 18650 -2200
rect 18730 -2240 18790 -2160
rect 18510 -2260 18790 -2240
rect 18510 -2320 18530 -2260
rect 18590 -2320 18790 -2260
rect 18510 -2350 18790 -2320
rect 2360 -3100 2760 -3080
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3340 2760 -3280
rect 2360 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect 2360 -3480 2760 -3420
rect -5170 -3760 -1570 -3560
rect -5170 -17300 -4770 -3760
rect -2320 -4220 -1920 -4190
rect -2320 -4300 -2290 -4220
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -2320 -4370 -1920 -4300
rect -2320 -4450 -2290 -4370
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -2320 -4490 -1920 -4450
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4590 -1920 -4550
rect -1770 -4210 -1570 -3760
rect 13160 -3570 13420 -3540
rect 13160 -3580 13300 -3570
rect 13160 -3640 13170 -3580
rect 13230 -3640 13300 -3580
rect 13160 -3650 13300 -3640
rect 13380 -3650 13420 -3570
rect 13160 -3700 13420 -3650
rect 13160 -3760 13170 -3700
rect 13230 -3760 13420 -3700
rect 13160 -3810 13420 -3760
rect 13160 -3890 13300 -3810
rect 13380 -3890 13420 -3810
rect 13160 -3940 13420 -3890
rect -1770 -4310 -1730 -4210
rect -1630 -4310 -1570 -4210
rect -1770 -4380 -1570 -4310
rect -1770 -4480 -1730 -4380
rect -1630 -4480 -1570 -4380
rect -1770 -4540 -1570 -4480
rect -1770 -4640 -1730 -4540
rect -1630 -4640 -1570 -4540
rect -1770 -4660 -1570 -4640
rect 4530 -4480 6740 -4460
rect 4530 -4540 6560 -4480
rect 6620 -4540 6660 -4480
rect 6720 -4540 6740 -4480
rect 4530 -4580 6740 -4540
rect 4530 -4640 6560 -4580
rect 6620 -4640 6660 -4580
rect 6720 -4640 6740 -4580
rect 4530 -4660 6740 -4640
rect -1480 -5500 -1080 -5470
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5630 -1080 -5560
rect -1480 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 -1080 -5630
rect -1480 -5770 -1080 -5710
rect -1480 -5850 -1430 -5770
rect -1350 -5850 -1230 -5770
rect -1150 -5850 -1080 -5770
rect -1480 -5870 -1080 -5850
rect -90 -5500 310 -5470
rect -90 -5560 -60 -5500
rect 0 -5560 60 -5500
rect 120 -5560 180 -5500
rect 240 -5560 310 -5500
rect -90 -5630 310 -5560
rect -90 -5710 -40 -5630
rect 40 -5710 160 -5630
rect 240 -5710 310 -5630
rect -90 -5770 310 -5710
rect -90 -5850 -40 -5770
rect 40 -5850 160 -5770
rect 240 -5850 310 -5770
rect -90 -5870 310 -5850
rect 1060 -5690 3230 -5670
rect 1060 -5750 1080 -5690
rect 1140 -5750 1200 -5690
rect 1260 -5750 3230 -5690
rect 1060 -5790 3230 -5750
rect 1060 -5850 1080 -5790
rect 1140 -5850 1200 -5790
rect 1260 -5850 3230 -5790
rect 1060 -5870 3230 -5850
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7210 -1480 -7150
rect -1960 -7290 -1930 -7210
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -1960 -7320 -1480 -7290
rect 580 -9160 980 -9140
rect 580 -9220 610 -9160
rect 670 -9220 730 -9160
rect 790 -9220 850 -9160
rect 910 -9220 980 -9160
rect 580 -9260 980 -9220
rect 580 -9340 610 -9260
rect 690 -9340 840 -9260
rect 920 -9340 980 -9260
rect 580 -9360 980 -9340
rect -3060 -9390 -2660 -9370
rect -3060 -9450 -3030 -9390
rect -2970 -9450 -2910 -9390
rect -2850 -9450 -2790 -9390
rect -2730 -9450 -2660 -9390
rect -3060 -9480 -2660 -9450
rect -3060 -9560 -3030 -9480
rect -2950 -9560 -2800 -9480
rect -2720 -9560 -2660 -9480
rect -3060 -9590 -2660 -9560
rect -5170 -17460 -3380 -17300
rect -5170 -17700 -3386 -17460
rect -7590 -18966 -7038 -17770
rect -3938 -18966 -3386 -17700
rect 2830 -17770 3230 -5870
rect 2806 -18966 3358 -17770
rect 4530 -63620 4930 -4660
rect 9100 -4890 11680 -4690
rect 9100 -4950 9300 -4890
rect 9100 -5010 9120 -4950
rect 9180 -5010 9220 -4950
rect 9280 -5010 9300 -4950
rect 9100 -5050 9300 -5010
rect 9100 -5110 9120 -5050
rect 9180 -5110 9220 -5050
rect 9280 -5110 9300 -5050
rect 9100 -5130 9300 -5110
rect 8000 -9580 8390 -9560
rect 8000 -9640 8030 -9580
rect 8090 -9640 8150 -9580
rect 8210 -9640 8270 -9580
rect 8330 -9640 8390 -9580
rect 8000 -9690 8390 -9640
rect 8000 -9770 8040 -9690
rect 8120 -9770 8260 -9690
rect 8340 -9770 8390 -9690
rect 8000 -9800 8390 -9770
rect 11480 -10560 11680 -4890
rect 18510 -7010 18760 -6940
rect 18510 -7070 18530 -7010
rect 18590 -7070 18760 -7010
rect 18510 -7130 18650 -7070
rect 18510 -7190 18530 -7130
rect 18590 -7150 18650 -7130
rect 18730 -7150 18760 -7070
rect 18590 -7190 18760 -7150
rect 18510 -7230 18760 -7190
rect 18510 -7250 18650 -7230
rect 18510 -7310 18530 -7250
rect 18590 -7310 18650 -7250
rect 18730 -7310 18760 -7230
rect 18510 -7340 18760 -7310
rect 12250 -8140 12650 -8120
rect 12250 -8200 12280 -8140
rect 12340 -8200 12400 -8140
rect 12460 -8200 12520 -8140
rect 12580 -8200 12650 -8140
rect 12250 -8230 12650 -8200
rect 12250 -8310 12270 -8230
rect 12350 -8310 12510 -8230
rect 12590 -8310 12650 -8230
rect 12250 -8320 12650 -8310
rect 16070 -9580 16460 -9560
rect 16070 -9640 16090 -9580
rect 16150 -9640 16210 -9580
rect 16270 -9640 16330 -9580
rect 16390 -9640 16460 -9580
rect 16070 -9690 16460 -9640
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9800 16460 -9770
rect 11480 -10650 26430 -10560
rect 11480 -10850 25080 -10650
rect 25280 -10850 25480 -10650
rect 25680 -10850 25880 -10650
rect 26080 -10850 26430 -10650
rect 11480 -10970 26430 -10850
rect 4530 -63720 26670 -63620
rect 4530 -63920 25350 -63720
rect 25550 -63920 25750 -63720
rect 25950 -63920 26150 -63720
rect 26350 -63920 26670 -63720
rect 4530 -64020 26670 -63920
<< via2 >>
rect -250 8100 -170 8180
rect -10 8100 70 8180
rect 3060 8110 3140 8190
rect 3280 8110 3360 8190
rect 11080 8110 11160 8190
rect 11310 8110 11390 8190
rect 15900 8100 15980 8180
rect 16140 8100 16220 8180
rect 14830 4470 14930 4570
rect 14830 4270 14930 4370
rect -1430 880 -1350 960
rect -1220 880 -1140 960
rect -1430 740 -1350 820
rect -1220 740 -1140 820
rect -270 870 -190 950
rect -50 870 30 950
rect -270 730 -190 810
rect -50 730 30 810
rect 930 900 1010 980
rect 1170 900 1250 980
rect 930 740 1010 820
rect 1170 740 1250 820
rect 18650 -2080 18730 -2000
rect 18650 -2240 18730 -2160
rect 2380 -3420 2460 -3340
rect 2540 -3420 2620 -3340
rect -2290 -4300 -2210 -4220
rect -2040 -4300 -1960 -4220
rect -2290 -4450 -2210 -4370
rect -2040 -4450 -1960 -4370
rect 13300 -3650 13380 -3570
rect 13300 -3890 13380 -3810
rect -1430 -5710 -1350 -5630
rect -1230 -5710 -1150 -5630
rect -1430 -5850 -1350 -5770
rect -1230 -5850 -1150 -5770
rect -40 -5710 40 -5630
rect 160 -5710 240 -5630
rect -40 -5850 40 -5770
rect 160 -5850 240 -5770
rect -1930 -7290 -1850 -7210
rect -1770 -7290 -1690 -7210
rect -1610 -7290 -1530 -7210
rect 610 -9340 690 -9260
rect 840 -9340 920 -9260
rect -3030 -9560 -2950 -9480
rect -2800 -9560 -2720 -9480
rect 8040 -9770 8120 -9690
rect 8260 -9770 8340 -9690
rect 18650 -7150 18730 -7070
rect 18650 -7310 18730 -7230
rect 12270 -8310 12350 -8230
rect 12510 -8310 12590 -8230
rect 16100 -9770 16180 -9690
rect 16340 -9770 16420 -9690
rect 25080 -10850 25280 -10650
rect 25480 -10850 25680 -10650
rect 25880 -10850 26080 -10650
rect 25350 -63920 25550 -63720
rect 25750 -63920 25950 -63720
rect 26150 -63920 26350 -63720
<< metal3 >>
rect -6324 11740 22920 11900
rect -6324 11640 -6240 11740
rect -6140 11640 -6040 11740
rect -5940 11730 15920 11740
rect -5940 11640 -250 11730
rect -6324 11630 -250 11640
rect -150 11630 -50 11730
rect 50 11630 3060 11730
rect 3160 11630 3260 11730
rect 3360 11630 11080 11730
rect 11180 11630 11280 11730
rect 11380 11640 15920 11730
rect 16020 11640 16120 11740
rect 16220 11730 22920 11740
rect 16220 11640 22440 11730
rect 11380 11630 22440 11640
rect 22540 11630 22640 11730
rect 22740 11630 22920 11730
rect -6324 11540 22920 11630
rect -6324 11440 -6240 11540
rect -6140 11440 -6040 11540
rect -5940 11530 15920 11540
rect -5940 11440 -250 11530
rect -6324 11430 -250 11440
rect -150 11430 -50 11530
rect 50 11430 3060 11530
rect 3160 11430 3260 11530
rect 3360 11430 11080 11530
rect 11180 11430 11280 11530
rect 11380 11440 15920 11530
rect 16020 11440 16120 11540
rect 16220 11530 22920 11540
rect 16220 11440 22440 11530
rect 11380 11430 22440 11440
rect 22540 11430 22640 11530
rect 22740 11430 22920 11530
rect -6324 11356 22920 11430
rect -4148 10300 21220 10420
rect -4148 10200 -4070 10300
rect -3970 10200 -3870 10300
rect -3770 10290 21220 10300
rect -3770 10200 20860 10290
rect -4148 10190 20860 10200
rect 20960 10190 21060 10290
rect 21160 10190 21220 10290
rect -4148 10100 21220 10190
rect -4148 10000 -4070 10100
rect -3970 10000 -3870 10100
rect -3770 10090 21220 10100
rect -3770 10000 20860 10090
rect -4148 9990 20860 10000
rect 20960 9990 21060 10090
rect 21160 9990 21220 10090
rect -4148 9876 21220 9990
rect 3020 8350 3420 8370
rect 3020 8250 3060 8350
rect 3160 8250 3260 8350
rect 3360 8250 3420 8350
rect -290 8200 110 8210
rect -290 8080 -270 8200
rect -150 8080 -30 8200
rect 90 8080 110 8200
rect -290 8070 110 8080
rect 3020 8190 3420 8250
rect 3020 8110 3060 8190
rect 3140 8110 3280 8190
rect 3360 8110 3420 8190
rect 3020 8070 3420 8110
rect 11040 8350 11440 8370
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 8190 11440 8250
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8070 11440 8110
rect 15870 8330 16270 8350
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 8180 16270 8230
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8070 16270 8100
rect 14680 4570 21210 4630
rect 14680 4470 14830 4570
rect 14930 4470 20760 4570
rect 20860 4470 21060 4570
rect 21160 4470 21210 4570
rect 14680 4370 21210 4470
rect 14680 4270 14830 4370
rect 14930 4270 20760 4370
rect 20860 4270 21060 4370
rect 21160 4270 21210 4370
rect 14680 4230 21210 4270
rect -6290 1050 1290 1110
rect -6290 950 -6250 1050
rect -6150 950 -6050 1050
rect -5950 980 1290 1050
rect -5950 960 930 980
rect -5950 950 -1430 960
rect -6290 880 -1430 950
rect -1350 880 -1220 960
rect -1140 950 930 960
rect -1140 880 -270 950
rect -6290 870 -270 880
rect -190 870 -50 950
rect 30 900 930 950
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 30 870 1290 900
rect -6290 850 1290 870
rect -6290 750 -6250 850
rect -6150 750 -6050 850
rect -5950 820 1290 850
rect -5950 750 -1430 820
rect -6290 740 -1430 750
rect -1350 740 -1220 820
rect -1140 810 930 820
rect -1140 740 -270 810
rect -6290 730 -270 740
rect -190 730 -50 810
rect 30 740 930 810
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 30 730 1290 740
rect -6290 710 1290 730
rect 18510 -2000 21210 -1950
rect 18510 -2080 18650 -2000
rect 18730 -2080 20870 -2000
rect 18510 -2100 20870 -2080
rect 20970 -2100 21070 -2000
rect 21170 -2100 21210 -2000
rect 18510 -2160 21210 -2100
rect 18510 -2240 18650 -2160
rect 18730 -2200 21210 -2160
rect 18730 -2240 20870 -2200
rect 18510 -2300 20870 -2240
rect 20970 -2300 21070 -2200
rect 21170 -2300 21210 -2200
rect 18510 -2350 21210 -2300
rect -4130 -3120 2760 -3080
rect -4130 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 2760 -3120
rect -4130 -3320 2760 -3220
rect -4130 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3340 2760 -3320
rect -3770 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect -4130 -3480 2760 -3420
rect 13160 -3570 22920 -3540
rect 13160 -3650 13300 -3570
rect 13380 -3580 22920 -3570
rect 13380 -3650 22450 -3580
rect 13160 -3680 22450 -3650
rect 22550 -3680 22650 -3580
rect 22750 -3680 22920 -3580
rect 13160 -3780 22920 -3680
rect 13160 -3810 22450 -3780
rect 13160 -3890 13300 -3810
rect 13380 -3880 22450 -3810
rect 22550 -3880 22650 -3780
rect 22750 -3880 22920 -3780
rect 13380 -3890 22920 -3880
rect 13160 -3940 22920 -3890
rect -6290 -4220 -1920 -4190
rect -6290 -4230 -2290 -4220
rect -6290 -4330 -6240 -4230
rect -6140 -4330 -6040 -4230
rect -5940 -4300 -2290 -4230
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -5940 -4330 -1920 -4300
rect -6290 -4370 -1920 -4330
rect -6290 -4430 -2290 -4370
rect -6290 -4530 -6240 -4430
rect -6140 -4530 -6040 -4430
rect -5940 -4450 -2290 -4430
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -5940 -4530 -1920 -4450
rect -6290 -4590 -1920 -4530
rect -4130 -5520 310 -5470
rect -4130 -5620 -4090 -5520
rect -3990 -5620 -3890 -5520
rect -3790 -5620 310 -5520
rect -4130 -5630 310 -5620
rect -4130 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 -40 -5630
rect 40 -5710 160 -5630
rect 240 -5710 310 -5630
rect -4130 -5720 310 -5710
rect -4130 -5820 -4090 -5720
rect -3990 -5820 -3890 -5720
rect -3790 -5770 310 -5720
rect -3790 -5820 -1430 -5770
rect -4130 -5850 -1430 -5820
rect -1350 -5850 -1230 -5770
rect -1150 -5850 -40 -5770
rect 40 -5850 160 -5770
rect 240 -5850 310 -5770
rect -4130 -5870 310 -5850
rect 18510 -6990 21210 -6940
rect -4130 -7080 -1480 -7030
rect -4130 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -1480 -7080
rect -4130 -7210 -1480 -7180
rect -4130 -7280 -1930 -7210
rect -4130 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7290 -1930 -7280
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -3790 -7320 -1480 -7290
rect 18510 -7070 20860 -6990
rect 18510 -7150 18650 -7070
rect 18730 -7090 20860 -7070
rect 20960 -7090 21060 -6990
rect 21160 -7090 21210 -6990
rect 18730 -7150 21210 -7090
rect 18510 -7190 21210 -7150
rect 18510 -7230 20860 -7190
rect 18510 -7310 18650 -7230
rect 18730 -7290 20860 -7230
rect 20960 -7290 21060 -7190
rect 21160 -7290 21210 -7190
rect 18730 -7310 21210 -7290
rect -3790 -7380 -3730 -7320
rect 18510 -7340 21210 -7310
rect -4130 -7430 -3730 -7380
rect 12250 -8230 12650 -8220
rect 12250 -8310 12270 -8230
rect 12350 -8310 12510 -8230
rect 12590 -8310 12650 -8230
rect 12250 -8330 12650 -8310
rect 12250 -8430 12280 -8330
rect 12380 -8430 12480 -8330
rect 12580 -8430 12650 -8330
rect 12250 -8440 12650 -8430
rect 580 -9260 980 -9240
rect 580 -9340 610 -9260
rect 690 -9340 840 -9260
rect 920 -9340 980 -9260
rect 580 -9370 980 -9340
rect -3060 -9480 -2660 -9460
rect 580 -9470 600 -9370
rect 700 -9470 800 -9370
rect 900 -9470 980 -9370
rect 580 -9480 980 -9470
rect -3060 -9560 -3030 -9480
rect -2950 -9560 -2800 -9480
rect -2720 -9560 -2660 -9480
rect -3060 -9600 -2660 -9560
rect -3060 -9700 -3030 -9600
rect -2930 -9700 -2830 -9600
rect -2730 -9700 -2660 -9600
rect -3060 -9720 -2660 -9700
rect 8000 -9690 8390 -9660
rect 8000 -9770 8040 -9690
rect 8120 -9770 8260 -9690
rect 8340 -9770 8390 -9690
rect 8000 -9800 8390 -9770
rect 8000 -9900 8030 -9800
rect 8130 -9900 8250 -9800
rect 8350 -9900 8390 -9800
rect 8000 -9910 8390 -9900
rect 16070 -9690 16460 -9660
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9820 16460 -9770
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -9940 16460 -9920
rect 24888 -10650 26520 -10404
rect 24888 -10850 25080 -10650
rect 25280 -10850 25480 -10650
rect 25680 -10850 25880 -10650
rect 26080 -10850 26520 -10650
rect 24888 -11084 26520 -10850
rect -4148 -11510 21220 -11356
rect -4148 -11610 -4070 -11510
rect -3970 -11610 -3870 -11510
rect -3770 -11520 21220 -11510
rect -3770 -11610 8040 -11520
rect -4148 -11620 8040 -11610
rect 8140 -11620 8240 -11520
rect 8340 -11620 16120 -11520
rect 16220 -11620 16320 -11520
rect 16420 -11530 21220 -11520
rect 16420 -11620 20850 -11530
rect -4148 -11630 20850 -11620
rect 20950 -11630 21050 -11530
rect 21150 -11630 21220 -11530
rect -4148 -11710 21220 -11630
rect -4148 -11810 -4070 -11710
rect -3970 -11810 -3870 -11710
rect -3770 -11720 21220 -11710
rect -3770 -11810 8040 -11720
rect -4148 -11820 8040 -11810
rect 8140 -11820 8240 -11720
rect 8340 -11820 16120 -11720
rect 16220 -11820 16320 -11720
rect 16420 -11730 21220 -11720
rect 16420 -11820 20850 -11730
rect -4148 -11830 20850 -11820
rect 20950 -11830 21050 -11730
rect 21150 -11830 21220 -11730
rect -4148 -11900 21220 -11830
rect -6324 -13710 22920 -13532
rect -6324 -13720 630 -13710
rect -6324 -13820 -6240 -13720
rect -6140 -13820 -6040 -13720
rect -5940 -13730 630 -13720
rect -5940 -13820 -3000 -13730
rect -6324 -13830 -3000 -13820
rect -2900 -13830 -2800 -13730
rect -2700 -13810 630 -13730
rect 730 -13810 830 -13710
rect 930 -13810 12300 -13710
rect 12400 -13810 12500 -13710
rect 12600 -13730 22920 -13710
rect 12600 -13810 22440 -13730
rect -2700 -13830 22440 -13810
rect 22540 -13830 22640 -13730
rect 22740 -13830 22920 -13730
rect -6324 -13910 22920 -13830
rect -6324 -13920 630 -13910
rect -6324 -14020 -6240 -13920
rect -6140 -14020 -6040 -13920
rect -5940 -13930 630 -13920
rect -5940 -14020 -3000 -13930
rect -6324 -14030 -3000 -14020
rect -2900 -14030 -2800 -13930
rect -2700 -14010 630 -13930
rect 730 -14010 830 -13910
rect 930 -14010 12300 -13910
rect 12400 -14010 12500 -13910
rect 12600 -13930 22920 -13910
rect 12600 -14010 22440 -13930
rect -2700 -14030 22440 -14010
rect 22540 -14030 22640 -13930
rect 22740 -14030 22920 -13930
rect -6324 -14076 22920 -14030
rect 25092 -63720 26724 -63580
rect 25092 -63920 25350 -63720
rect 25550 -63920 25750 -63720
rect 25950 -63920 26150 -63720
rect 26350 -63920 26724 -63720
rect 25092 -64124 26724 -63920
<< via3 >>
rect -6240 11640 -6140 11740
rect -6040 11640 -5940 11740
rect -250 11630 -150 11730
rect -50 11630 50 11730
rect 3060 11630 3160 11730
rect 3260 11630 3360 11730
rect 11080 11630 11180 11730
rect 11280 11630 11380 11730
rect 15920 11640 16020 11740
rect 16120 11640 16220 11740
rect 22440 11630 22540 11730
rect 22640 11630 22740 11730
rect -6240 11440 -6140 11540
rect -6040 11440 -5940 11540
rect -250 11430 -150 11530
rect -50 11430 50 11530
rect 3060 11430 3160 11530
rect 3260 11430 3360 11530
rect 11080 11430 11180 11530
rect 11280 11430 11380 11530
rect 15920 11440 16020 11540
rect 16120 11440 16220 11540
rect 22440 11430 22540 11530
rect 22640 11430 22740 11530
rect -4070 10200 -3970 10300
rect -3870 10200 -3770 10300
rect 20860 10190 20960 10290
rect 21060 10190 21160 10290
rect -4070 10000 -3970 10100
rect -3870 10000 -3770 10100
rect 20860 9990 20960 10090
rect 21060 9990 21160 10090
rect 3060 8250 3160 8350
rect 3260 8250 3360 8350
rect -270 8180 -150 8200
rect -270 8100 -250 8180
rect -250 8100 -170 8180
rect -170 8100 -150 8180
rect -270 8080 -150 8100
rect -30 8180 90 8200
rect -30 8100 -10 8180
rect -10 8100 70 8180
rect 70 8100 90 8180
rect -30 8080 90 8100
rect 11080 8250 11180 8350
rect 11280 8250 11380 8350
rect 15900 8230 16000 8330
rect 16130 8230 16230 8330
rect 20760 4470 20860 4570
rect 21060 4470 21160 4570
rect 20760 4270 20860 4370
rect 21060 4270 21160 4370
rect -6250 950 -6150 1050
rect -6050 950 -5950 1050
rect -6250 750 -6150 850
rect -6050 750 -5950 850
rect 20870 -2100 20970 -2000
rect 21070 -2100 21170 -2000
rect 20870 -2300 20970 -2200
rect 21070 -2300 21170 -2200
rect -4070 -3220 -3970 -3120
rect -3870 -3220 -3770 -3120
rect -4070 -3420 -3970 -3320
rect -3870 -3420 -3770 -3320
rect 22450 -3680 22550 -3580
rect 22650 -3680 22750 -3580
rect 22450 -3880 22550 -3780
rect 22650 -3880 22750 -3780
rect -6240 -4330 -6140 -4230
rect -6040 -4330 -5940 -4230
rect -6240 -4530 -6140 -4430
rect -6040 -4530 -5940 -4430
rect -4090 -5620 -3990 -5520
rect -3890 -5620 -3790 -5520
rect -4090 -5820 -3990 -5720
rect -3890 -5820 -3790 -5720
rect -4090 -7180 -3990 -7080
rect -3890 -7180 -3790 -7080
rect -4090 -7380 -3990 -7280
rect -3890 -7380 -3790 -7280
rect 20860 -7090 20960 -6990
rect 21060 -7090 21160 -6990
rect 20860 -7290 20960 -7190
rect 21060 -7290 21160 -7190
rect 12280 -8430 12380 -8330
rect 12480 -8430 12580 -8330
rect 600 -9470 700 -9370
rect 800 -9470 900 -9370
rect -3030 -9700 -2930 -9600
rect -2830 -9700 -2730 -9600
rect 8030 -9900 8130 -9800
rect 8250 -9900 8350 -9800
rect 16110 -9920 16210 -9820
rect 16310 -9920 16410 -9820
rect -4070 -11610 -3970 -11510
rect -3870 -11610 -3770 -11510
rect 8040 -11620 8140 -11520
rect 8240 -11620 8340 -11520
rect 16120 -11620 16220 -11520
rect 16320 -11620 16420 -11520
rect 20850 -11630 20950 -11530
rect 21050 -11630 21150 -11530
rect -4070 -11810 -3970 -11710
rect -3870 -11810 -3770 -11710
rect 8040 -11820 8140 -11720
rect 8240 -11820 8340 -11720
rect 16120 -11820 16220 -11720
rect 16320 -11820 16420 -11720
rect 20850 -11830 20950 -11730
rect 21050 -11830 21150 -11730
rect -6240 -13820 -6140 -13720
rect -6040 -13820 -5940 -13720
rect -3000 -13830 -2900 -13730
rect -2800 -13830 -2700 -13730
rect 630 -13810 730 -13710
rect 830 -13810 930 -13710
rect 12300 -13810 12400 -13710
rect 12500 -13810 12600 -13710
rect 22440 -13830 22540 -13730
rect 22640 -13830 22740 -13730
rect -6240 -14020 -6140 -13920
rect -6040 -14020 -5940 -13920
rect -3000 -14030 -2900 -13930
rect -2800 -14030 -2700 -13930
rect 630 -14010 730 -13910
rect 830 -14010 930 -13910
rect 12300 -14010 12400 -13910
rect 12500 -14010 12600 -13910
rect 22440 -14030 22540 -13930
rect 22640 -14030 22740 -13930
<< metal4 >>
rect -6324 11740 -5780 11900
rect -6324 11640 -6240 11740
rect -6140 11640 -6040 11740
rect -5940 11640 -5780 11740
rect -6324 11540 -5780 11640
rect -6324 11440 -6240 11540
rect -6140 11440 -6040 11540
rect -5940 11440 -5780 11540
rect -6324 1050 -5780 11440
rect -300 11790 100 11900
rect -300 11730 110 11790
rect -300 11630 -250 11730
rect -150 11630 -50 11730
rect 50 11630 110 11730
rect -300 11530 110 11630
rect -300 11430 -250 11530
rect -150 11430 -50 11530
rect 50 11430 110 11530
rect -300 11340 110 11430
rect 3020 11730 3420 11790
rect 3020 11630 3060 11730
rect 3160 11630 3260 11730
rect 3360 11630 3420 11730
rect 3020 11530 3420 11630
rect 3020 11430 3060 11530
rect 3160 11430 3260 11530
rect 3360 11430 3420 11530
rect -6324 950 -6250 1050
rect -6150 950 -6050 1050
rect -5950 950 -5780 1050
rect -6324 850 -5780 950
rect -6324 750 -6250 850
rect -6150 750 -6050 850
rect -5950 750 -5780 850
rect -6324 -4230 -5780 750
rect -6324 -4330 -6240 -4230
rect -6140 -4330 -6040 -4230
rect -5940 -4330 -5780 -4230
rect -6324 -4430 -5780 -4330
rect -6324 -4530 -6240 -4430
rect -6140 -4530 -6040 -4430
rect -5940 -4530 -5780 -4430
rect -6324 -13720 -5780 -4530
rect -4148 10300 -3604 10420
rect -4148 10200 -4070 10300
rect -3970 10200 -3870 10300
rect -3770 10200 -3604 10300
rect -4148 10100 -3604 10200
rect -4148 10000 -4070 10100
rect -3970 10000 -3870 10100
rect -3770 10000 -3604 10100
rect -4148 -3120 -3604 10000
rect -300 8260 100 11340
rect 3020 8350 3420 11430
rect -300 8240 110 8260
rect -290 8200 110 8240
rect -290 8080 -270 8200
rect -150 8080 -30 8200
rect 90 8080 110 8200
rect -290 7990 110 8080
rect 3020 8250 3060 8350
rect 3160 8250 3260 8350
rect 3360 8250 3420 8350
rect 3020 7990 3420 8250
rect 11040 11730 11440 11790
rect 11040 11630 11080 11730
rect 11180 11630 11280 11730
rect 11380 11630 11440 11730
rect 11040 11530 11440 11630
rect 11040 11430 11080 11530
rect 11180 11430 11280 11530
rect 11380 11430 11440 11530
rect 11040 8350 11440 11430
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 7990 11440 8250
rect 15870 11740 16270 11790
rect 15870 11640 15920 11740
rect 16020 11640 16120 11740
rect 16220 11640 16270 11740
rect 15870 11540 16270 11640
rect 15870 11440 15920 11540
rect 16020 11440 16120 11540
rect 16220 11440 16270 11540
rect 15870 8330 16270 11440
rect 22376 11730 22920 11900
rect 22376 11630 22440 11730
rect 22540 11630 22640 11730
rect 22740 11630 22920 11730
rect 22376 11530 22920 11630
rect 22376 11430 22440 11530
rect 22540 11430 22640 11530
rect 22740 11430 22920 11530
rect 22376 11340 22920 11430
rect 20676 10290 21220 10420
rect 20676 10190 20860 10290
rect 20960 10190 21060 10290
rect 21160 10190 21220 10290
rect 20676 10090 21220 10190
rect 20676 9990 20860 10090
rect 20960 9990 21060 10090
rect 21160 9990 21220 10090
rect 20676 9860 21220 9990
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 7990 16270 8230
rect 20680 4640 21220 9860
rect 20676 4570 21220 4640
rect 20676 4470 20760 4570
rect 20860 4470 21060 4570
rect 21160 4470 21220 4570
rect 20676 4370 21220 4470
rect 20676 4270 20760 4370
rect 20860 4270 21060 4370
rect 21160 4270 21220 4370
rect 20676 4220 21220 4270
rect 20680 -1940 21220 4220
rect 20676 -2000 21220 -1940
rect 20676 -2100 20870 -2000
rect 20970 -2100 21070 -2000
rect 21170 -2100 21220 -2000
rect 20676 -2200 21220 -2100
rect 20676 -2300 20870 -2200
rect 20970 -2300 21070 -2200
rect 21170 -2300 21220 -2200
rect 20676 -2360 21220 -2300
rect -4148 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 -3604 -3120
rect -4148 -3320 -3604 -3220
rect -4148 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3420 -3604 -3320
rect -4148 -5520 -3604 -3420
rect -4148 -5620 -4090 -5520
rect -3990 -5620 -3890 -5520
rect -3790 -5620 -3604 -5520
rect -4148 -5720 -3604 -5620
rect -4148 -5820 -4090 -5720
rect -3990 -5820 -3890 -5720
rect -3790 -5820 -3604 -5720
rect -4148 -7080 -3604 -5820
rect 20680 -6940 21220 -2360
rect 22380 -3540 22920 11340
rect 22376 -3580 22920 -3540
rect 22376 -3680 22450 -3580
rect 22550 -3680 22650 -3580
rect 22750 -3680 22920 -3580
rect 22376 -3780 22920 -3680
rect 22376 -3880 22450 -3780
rect 22550 -3880 22650 -3780
rect 22750 -3880 22920 -3780
rect 22376 -3940 22920 -3880
rect -4148 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -3604 -7080
rect -4148 -7280 -3604 -7180
rect -4148 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7380 -3604 -7280
rect 20676 -6990 21220 -6940
rect 20676 -7090 20860 -6990
rect 20960 -7090 21060 -6990
rect 21160 -7090 21220 -6990
rect 20676 -7190 21220 -7090
rect 20676 -7290 20860 -7190
rect 20960 -7290 21060 -7190
rect 21160 -7290 21220 -7190
rect 20676 -7340 21220 -7290
rect -4148 -11510 -3604 -7380
rect 12250 -8330 12650 -8120
rect 12250 -8430 12280 -8330
rect 12380 -8430 12480 -8330
rect 12580 -8430 12650 -8330
rect 580 -9370 980 -9140
rect -4148 -11610 -4070 -11510
rect -3970 -11610 -3870 -11510
rect -3770 -11610 -3604 -11510
rect -4148 -11710 -3604 -11610
rect -4148 -11810 -4070 -11710
rect -3970 -11810 -3870 -11710
rect -3770 -11810 -3604 -11710
rect -4148 -11900 -3604 -11810
rect -3060 -9600 -2660 -9370
rect -3060 -9700 -3030 -9600
rect -2930 -9700 -2830 -9600
rect -2730 -9700 -2660 -9600
rect 580 -9470 600 -9370
rect 700 -9470 800 -9370
rect 900 -9470 980 -9370
rect -6324 -13820 -6240 -13720
rect -6140 -13820 -6040 -13720
rect -5940 -13820 -5780 -13720
rect -6324 -13920 -5780 -13820
rect -6324 -14020 -6240 -13920
rect -6140 -14020 -6040 -13920
rect -5940 -14020 -5780 -13920
rect -6324 -14076 -5780 -14020
rect -3060 -13730 -2640 -9700
rect -3060 -13830 -3000 -13730
rect -2900 -13830 -2800 -13730
rect -2700 -13830 -2640 -13730
rect -3060 -13930 -2640 -13830
rect -3060 -14030 -3000 -13930
rect -2900 -14030 -2800 -13930
rect -2700 -14030 -2640 -13930
rect -3060 -14080 -2640 -14030
rect 580 -13710 980 -9470
rect 8000 -9800 8390 -9550
rect 8000 -9900 8030 -9800
rect 8130 -9900 8250 -9800
rect 8350 -9900 8390 -9800
rect 8000 -11520 8390 -9900
rect 8000 -11620 8040 -11520
rect 8140 -11620 8240 -11520
rect 8340 -11620 8390 -11520
rect 8000 -11720 8390 -11620
rect 8000 -11820 8040 -11720
rect 8140 -11820 8240 -11720
rect 8340 -11820 8390 -11720
rect 8000 -11870 8390 -11820
rect 580 -13810 630 -13710
rect 730 -13810 830 -13710
rect 930 -13810 980 -13710
rect 580 -13910 980 -13810
rect 580 -14010 630 -13910
rect 730 -14010 830 -13910
rect 930 -14010 980 -13910
rect 580 -14070 980 -14010
rect 12250 -13710 12650 -8430
rect 16070 -9820 16460 -9560
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -11520 16460 -9920
rect 20680 -11340 21220 -7340
rect 16070 -11620 16120 -11520
rect 16220 -11620 16320 -11520
rect 16420 -11620 16460 -11520
rect 16070 -11720 16460 -11620
rect 16070 -11820 16120 -11720
rect 16220 -11820 16320 -11720
rect 16420 -11820 16460 -11720
rect 16070 -11870 16460 -11820
rect 20676 -11530 21220 -11340
rect 20676 -11630 20850 -11530
rect 20950 -11630 21050 -11530
rect 21150 -11630 21220 -11530
rect 20676 -11730 21220 -11630
rect 20676 -11830 20850 -11730
rect 20950 -11830 21050 -11730
rect 21150 -11830 21220 -11730
rect 20676 -11900 21220 -11830
rect 22380 -13520 22920 -3940
rect 12250 -13810 12300 -13710
rect 12400 -13810 12500 -13710
rect 12600 -13810 12650 -13710
rect 12250 -13910 12650 -13810
rect 12250 -14010 12300 -13910
rect 12400 -14010 12500 -13910
rect 12600 -14010 12650 -13910
rect 12250 -14070 12650 -14010
rect 22376 -13730 22920 -13520
rect 22376 -13830 22440 -13730
rect 22540 -13830 22640 -13730
rect 22740 -13830 22920 -13730
rect 22376 -13930 22920 -13830
rect 22376 -14030 22440 -13930
rect 22540 -14030 22640 -13930
rect 22740 -14030 22920 -13930
rect 22376 -14076 22920 -14030
use ALib_DCO  ALib_DCO_0 ./../dco
timestamp 1730531556
transform 1 0 5200 0 1 -5190
box 1000 -4470 13410 5980
use ALib_VCO  ALib_VCO_0 ./../vco
timestamp 1730639796
transform 1 0 -2020 0 1 1040
box 0 280 20640 7030
use DLib_Quantizer  DLib_Quantizer_0 ./../quantizer
timestamp 1730532965
transform 1 0 -2210 0 1 -4630
box 190 -710 5890 730
use DLib_UpDownCounter  DLib_UpDownCounter_0 ./../count
timestamp 1730536752
transform 1 0 -1140 0 1 -5986
box -880 -3154 3140 -440
use DLib_UpDownCounter  DLib_UpDownCounter_1
timestamp 1730536752
transform 1 0 -1140 0 1 344
box -880 -3154 3140 -440
<< labels >>
flabel metal3 -5940 11356 -1070 11900 1 FreeSans 2176 0 0 0 VDDA
port 7 nsew power input
flabel metal3 25092 -64124 26724 -63580 1 FreeSans 1088 0 0 0 Vbs_12
port 1 nsew signal input
flabel metal2 17342 34914 17710 36938 1 FreeSans 736 0 0 0 Anlg_in
port 3 nsew signal input
flabel metal3 24888 -11084 26520 -10404 1 FreeSans 1088 0 0 0 Vbs_34
port 2 nsew signal input
flabel metal3 16388 9876 19516 10420 1 FreeSans 2176 0 0 0 GND
port 8 nsew ground input
flabel metal2 -7590 -18966 -7038 -17770 1 FreeSans 736 0 0 0 ENB
port 4 nsew signal input
flabel metal2 2806 -18966 3358 -17770 1 FreeSans 736 0 0 0 Dout
port 6 nsew signal input
flabel metal2 -3938 -18966 -3386 -17770 1 FreeSans 736 0 0 0 CLK
port 5 nsew signal input
<< end >>
