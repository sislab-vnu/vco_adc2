* this file contains all analog circuits written by SPICE

