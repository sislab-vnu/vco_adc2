* NGSPICE file created from p_br1.ext - technology: sky130A

.subckt p_br1 G S D B
X0 D G S B sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
.ends

