* NGSPICE file created from ALib_VCO.ext - technology: sky130A

.subckt aux_inv A Y VGND VDDA GND
X0 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt main_inv A Y VGND GND VDDA
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt cc_inv inp inn outp outn VGND GND VDDA
Xaux_inv_0 outp outn VGND VDDA GND aux_inv
Xaux_inv_1 outn outp VGND VDDA GND aux_inv
Xmain_inv_0 inp outp VGND GND VDDA main_inv
Xmain_inv_1 inn outn VGND GND VDDA main_inv
.ends

.subckt x5s_cc_osc pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VGND VDDA
+ GND
Xcc_inv_0 p[4] pn[4] p[0] pn[0] VGND GND VDDA cc_inv
Xcc_inv_1 p[0] pn[0] p[1] pn[1] VGND GND VDDA cc_inv
Xcc_inv_2 p[1] pn[1] p[2] pn[2] VGND GND VDDA cc_inv
Xcc_inv_3 p[3] pn[3] p[4] pn[4] VGND GND VDDA cc_inv
Xcc_inv_4 p[2] pn[2] p[3] pn[3] VGND GND VDDA cc_inv
.ends

.subckt sky130_fd_pr__res_generic_po_DKCPUZ a_n48_200# a_n48_n630#
R0 a_n48_200# a_n48_n630# sky130_fd_pr__res_generic_po w=0.48 l=2
.ends


.subckt ALib_VCO Anlg_in ENB p[4] VDDA GND
Xx5s_cc_osc_0 x5s_cc_osc_0/pn[0] x5s_cc_osc_0/pn[1] x5s_cc_osc_0/pn[2] x5s_cc_osc_0/pn[3]
+ pn[4] x5s_cc_osc_0/p[0] x5s_cc_osc_0/p[1] x5s_cc_osc_0/p[2] x5s_cc_osc_0/p[3] p[4]
+ Vctrl VDDA GND x5s_cc_osc
Xsky130_fd_pr__res_generic_po_DKCPUZ_0 Anlg_in Vctrl sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_pr__res_generic_po_DKCPUZ_1 Vctrl GND sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_sc_hd__einvp_1_0 VDDA ENB GND GND VDDA VDDA pn[4] sky130_fd_sc_hd__einvp_1
.ends


