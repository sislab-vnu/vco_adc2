magic
tech sky130A
timestamp 1725437652
<< nwell >>
rect 845 1055 865 1075
rect 2820 1055 2840 1075
rect 3710 1055 3730 1075
rect 5685 1055 5705 1075
rect 8550 1055 8570 1075
rect 845 1015 865 1035
rect 2820 1015 2840 1035
rect 5685 1015 5705 1035
rect 8550 1015 8570 1035
rect 2820 975 2840 995
rect 3710 975 3730 995
rect 835 965 875 970
rect 1840 -1605 1860 -1585
rect 3815 -1605 3835 -1585
rect 4705 -1605 4725 -1585
rect 6680 -1605 6700 -1585
rect 1840 -1645 1860 -1625
rect 3815 -1645 3835 -1625
rect 4705 -1645 4725 -1625
rect 6680 -1645 6700 -1625
rect 3815 -1685 3835 -1665
rect 4705 -1685 4725 -1665
rect 6680 -1685 6700 -1665
<< pwell >>
rect 845 170 865 190
rect 2820 170 2840 190
rect 3710 170 3730 190
rect 5685 170 5705 190
rect 6575 170 6595 190
rect 8550 170 8570 190
rect 845 130 865 150
rect 2820 130 2840 150
rect 3710 130 3730 150
rect 5685 130 5705 150
rect 6575 130 6595 150
rect 8550 130 8570 150
rect 845 90 865 110
rect 2820 90 2840 110
rect 20 20 105 85
rect 2880 20 2955 100
rect 5685 90 5705 110
rect 6575 90 6595 110
rect 5745 20 5805 65
rect 4605 -655 4670 -630
rect 7435 -680 7530 -630
rect 1840 -720 1860 -700
rect 3815 -720 3835 -700
rect 4705 -720 4725 -700
rect 6680 -720 6700 -700
rect 1840 -760 1860 -740
rect 3815 -760 3835 -740
rect 4705 -760 4725 -740
rect 6680 -760 6700 -740
rect 3815 -800 3835 -780
<< pdiff >>
rect 835 965 875 970
<< ndiffc >>
rect 845 170 865 190
rect 2820 170 2840 190
rect 3710 170 3730 190
rect 5685 170 5705 190
rect 6575 170 6595 190
rect 8550 170 8570 190
rect 845 130 865 150
rect 2820 130 2840 150
rect 3710 130 3730 150
rect 5685 130 5705 150
rect 6575 130 6595 150
rect 8550 130 8570 150
rect 845 90 865 110
rect 2820 90 2840 110
rect 5685 90 5705 110
rect 6575 90 6595 110
rect 1840 -720 1860 -700
rect 3815 -720 3835 -700
rect 4705 -720 4725 -700
rect 6680 -720 6700 -700
rect 1840 -760 1860 -740
rect 3815 -760 3835 -740
rect 4705 -760 4725 -740
rect 6680 -760 6700 -740
rect 3815 -800 3835 -780
<< pdiffc >>
rect 845 1055 865 1075
rect 2820 1055 2840 1075
rect 3710 1055 3730 1075
rect 5685 1055 5705 1075
rect 8550 1055 8570 1075
rect 845 1015 865 1035
rect 2820 1015 2840 1035
rect 5685 1015 5705 1035
rect 8550 1015 8570 1035
rect 2820 975 2840 995
rect 3710 975 3730 995
rect 1840 -1605 1860 -1585
rect 3815 -1605 3835 -1585
rect 4705 -1605 4725 -1585
rect 6680 -1605 6700 -1585
rect 1840 -1645 1860 -1625
rect 3815 -1645 3835 -1625
rect 4705 -1645 4725 -1625
rect 6680 -1645 6700 -1625
rect 3815 -1685 3835 -1665
rect 4705 -1685 4725 -1665
rect 6680 -1685 6700 -1665
<< locali >>
rect 80 1175 200 1215
rect 2825 1175 2910 1215
rect 5665 1175 5790 1215
rect 7630 1175 8580 1215
rect 905 1075 945 1090
rect 1930 1085 1970 1100
rect 3770 1075 3810 1090
rect 4795 1085 4835 1100
rect 6635 1075 6675 1090
rect 7660 1085 7700 1100
rect 835 965 875 970
rect 3770 80 3810 90
rect 4795 85 4835 90
rect 6635 80 6675 85
rect 905 45 945 80
rect 1830 -635 1870 -20
rect 2825 -50 2935 -10
rect 4615 -560 4655 -25
rect 5695 -50 5800 -10
rect 4585 -600 4750 -560
rect 4615 -635 4655 -600
rect 7480 -630 7520 -20
rect 2710 -695 2750 -690
rect 6600 -695 6640 -690
rect 2710 -1710 2750 -1695
rect 3735 -1700 3775 -1695
rect 1830 -1825 1905 -1785
rect 4640 -1825 4735 -1785
rect 7345 -1825 7520 -1785
<< viali >>
rect 845 1055 865 1075
rect 2820 1055 2840 1075
rect 3710 1055 3730 1075
rect 5685 1055 5705 1075
rect 8550 1055 8570 1075
rect 845 1015 865 1035
rect 2820 1015 2840 1035
rect 3710 1015 3730 1035
rect 5685 1015 5705 1035
rect 8550 1015 8570 1035
rect 845 975 865 995
rect 2820 975 2840 995
rect 3710 975 3730 995
rect 5685 975 5705 995
rect 8550 975 8570 995
rect 845 170 865 190
rect 2820 170 2840 190
rect 3710 170 3730 190
rect 5685 170 5705 190
rect 6575 170 6595 190
rect 8550 170 8570 190
rect 845 130 865 150
rect 2820 130 2840 150
rect 3710 130 3730 150
rect 5685 130 5705 150
rect 6575 130 6595 150
rect 8550 130 8570 150
rect 845 90 865 110
rect 2820 90 2840 110
rect 3710 90 3730 110
rect 5685 90 5705 110
rect 6575 90 6595 110
rect 8550 90 8570 110
rect 1840 -720 1860 -700
rect 3815 -720 3835 -700
rect 4705 -720 4725 -700
rect 6680 -720 6700 -700
rect 1840 -760 1860 -740
rect 3815 -760 3835 -740
rect 4705 -760 4725 -740
rect 6680 -760 6700 -740
rect 1840 -800 1860 -780
rect 3815 -800 3835 -780
rect 4705 -800 4725 -780
rect 6680 -800 6700 -780
rect 1840 -1605 1860 -1585
rect 3815 -1605 3835 -1585
rect 4705 -1605 4725 -1585
rect 6680 -1605 6700 -1585
rect 1840 -1645 1860 -1625
rect 3815 -1645 3835 -1625
rect 4705 -1645 4725 -1625
rect 6680 -1645 6700 -1625
rect 1840 -1685 1860 -1665
rect 3815 -1685 3835 -1665
rect 4705 -1685 4725 -1665
rect 6680 -1685 6700 -1665
<< metal1 >>
rect -705 1175 945 1230
rect -705 -1770 -650 1175
rect 905 1165 945 1175
rect 1930 1165 1970 1195
rect 835 1075 875 1085
rect 835 1055 845 1075
rect 865 1055 875 1075
rect 835 1035 875 1055
rect 835 1015 845 1035
rect 865 1015 875 1035
rect 835 995 875 1015
rect 835 975 845 995
rect 865 975 875 995
rect 835 965 875 975
rect 2810 1075 2850 1195
rect 3770 1090 3810 1195
rect 4795 1150 4835 1195
rect 6635 1165 6675 1195
rect 8540 1170 9305 1220
rect 2810 1055 2820 1075
rect 2840 1055 2850 1075
rect 2810 1035 2850 1055
rect 2810 1015 2820 1035
rect 2840 1015 2850 1035
rect 2810 995 2850 1015
rect 2810 975 2820 995
rect 2840 975 2850 995
rect 2810 965 2850 975
rect 3700 1075 3740 1085
rect 3700 1055 3710 1075
rect 3730 1055 3740 1075
rect 3700 1035 3740 1055
rect 3700 1015 3710 1035
rect 3730 1015 3740 1035
rect 3700 995 3740 1015
rect 3700 975 3710 995
rect 3730 975 3740 995
rect 3700 965 3740 975
rect 5675 1075 5715 1085
rect 5675 1055 5685 1075
rect 5705 1055 5715 1075
rect 5675 1035 5715 1055
rect 5675 1015 5685 1035
rect 5705 1015 5715 1035
rect 5675 995 5715 1015
rect 5675 975 5685 995
rect 5705 975 5715 995
rect 5675 965 5715 975
rect 8540 1075 8580 1170
rect 8540 1055 8550 1075
rect 8570 1055 8580 1075
rect 8540 1035 8580 1055
rect 8540 1015 8550 1035
rect 8570 1015 8580 1035
rect 8540 995 8580 1015
rect 8540 975 8550 995
rect 8570 975 8580 995
rect 8540 965 8580 975
rect -450 805 5 855
rect 8600 805 9055 855
rect -450 -1415 -395 805
rect -195 280 5 330
rect 8600 280 8805 330
rect -195 -890 -145 280
rect 835 190 875 200
rect 835 170 845 190
rect 865 170 875 190
rect 835 150 875 170
rect 835 130 845 150
rect 865 130 875 150
rect 835 110 875 130
rect 835 90 845 110
rect 865 90 875 110
rect 835 80 875 90
rect 2810 190 2850 200
rect 2810 170 2820 190
rect 2840 170 2850 190
rect 2810 150 2850 170
rect 2810 130 2820 150
rect 2840 130 2850 150
rect 2810 110 2850 130
rect 2810 90 2820 110
rect 2840 90 2850 110
rect 2810 80 2850 90
rect 3700 190 3740 200
rect 3700 170 3710 190
rect 3730 170 3740 190
rect 3700 150 3740 170
rect 3700 130 3710 150
rect 3730 130 3740 150
rect 3700 110 3740 130
rect 3700 90 3710 110
rect 3730 90 3740 110
rect 3700 80 3740 90
rect 5675 190 5715 200
rect 5675 170 5685 190
rect 5705 170 5715 190
rect 5675 150 5715 170
rect 5675 130 5685 150
rect 5705 130 5715 150
rect 5675 110 5715 130
rect 5675 90 5685 110
rect 5705 90 5715 110
rect 5675 80 5715 90
rect 6565 190 6605 200
rect 6565 170 6575 190
rect 6595 170 6605 190
rect 6565 150 6605 170
rect 6565 130 6575 150
rect 6595 130 6605 150
rect 6565 110 6605 130
rect 6565 90 6575 110
rect 6595 90 6605 110
rect 6565 80 6605 90
rect 8540 190 8580 200
rect 8540 170 8550 190
rect 8570 170 8580 190
rect 8540 150 8580 170
rect 8540 130 8550 150
rect 8570 130 8580 150
rect 8540 110 8580 130
rect 8540 90 8550 110
rect 8570 90 8580 110
rect 8540 80 8580 90
rect 905 -325 945 40
rect 1930 -325 1970 10
rect 3770 -325 3810 40
rect 4795 -325 4835 35
rect 6635 -325 6675 20
rect 7660 -325 7700 35
rect 905 -375 7700 -325
rect 2710 -655 2750 -375
rect 3735 -650 3775 -375
rect 5575 -635 5615 -375
rect 6600 -650 6640 -375
rect 1830 -700 1870 -690
rect 1830 -720 1840 -700
rect 1860 -720 1870 -700
rect 1830 -740 1870 -720
rect 1830 -760 1840 -740
rect 1860 -760 1870 -740
rect 1830 -780 1870 -760
rect 1830 -800 1840 -780
rect 1860 -800 1870 -780
rect 1830 -810 1870 -800
rect 3805 -700 3845 -690
rect 3805 -720 3815 -700
rect 3835 -720 3845 -700
rect 3805 -740 3845 -720
rect 3805 -760 3815 -740
rect 3835 -760 3845 -740
rect 3805 -780 3845 -760
rect 3805 -800 3815 -780
rect 3835 -800 3845 -780
rect 3805 -810 3845 -800
rect 4695 -700 4735 -690
rect 4695 -720 4705 -700
rect 4725 -720 4735 -700
rect 4695 -740 4735 -720
rect 4695 -760 4705 -740
rect 4725 -760 4735 -740
rect 4695 -780 4735 -760
rect 4695 -800 4705 -780
rect 4725 -800 4735 -780
rect 4695 -810 4735 -800
rect 6670 -700 6710 -690
rect 6670 -720 6680 -700
rect 6700 -720 6710 -700
rect 6670 -740 6710 -720
rect 6670 -760 6680 -740
rect 6700 -760 6710 -740
rect 6670 -780 6710 -760
rect 6670 -800 6680 -780
rect 6700 -800 6710 -780
rect 6670 -810 6710 -800
rect 8755 -890 8805 280
rect -195 -940 1810 -890
rect 7540 -940 8805 -890
rect 9005 -1415 9055 805
rect -450 -1465 1810 -1415
rect 7535 -1465 9055 -1415
rect 1830 -1585 1870 -1575
rect 1830 -1605 1840 -1585
rect 1860 -1605 1870 -1585
rect 1830 -1625 1870 -1605
rect 1830 -1645 1840 -1625
rect 1860 -1645 1870 -1625
rect 1830 -1665 1870 -1645
rect 1830 -1685 1840 -1665
rect 1860 -1685 1870 -1665
rect 1830 -1770 1870 -1685
rect 3805 -1585 3845 -1575
rect 3805 -1605 3815 -1585
rect 3835 -1605 3845 -1585
rect 3805 -1625 3845 -1605
rect 3805 -1645 3815 -1625
rect 3835 -1645 3845 -1625
rect 3805 -1665 3845 -1645
rect 3805 -1685 3815 -1665
rect 3835 -1685 3845 -1665
rect 3805 -1695 3845 -1685
rect 4695 -1585 4735 -1575
rect 4695 -1605 4705 -1585
rect 4725 -1605 4735 -1585
rect 4695 -1625 4735 -1605
rect 4695 -1645 4705 -1625
rect 4725 -1645 4735 -1625
rect 4695 -1665 4735 -1645
rect 4695 -1685 4705 -1665
rect 4725 -1685 4735 -1665
rect 4695 -1695 4735 -1685
rect 6670 -1585 6710 -1575
rect 6670 -1605 6680 -1585
rect 6700 -1605 6710 -1585
rect 6670 -1625 6710 -1605
rect 6670 -1645 6680 -1625
rect 6700 -1645 6710 -1625
rect 6670 -1665 6710 -1645
rect 6670 -1685 6680 -1665
rect 6700 -1685 6710 -1665
rect 6670 -1695 6710 -1685
rect -705 -1825 1870 -1770
rect 6600 -1775 6640 -1765
rect 9255 -1775 9305 1170
rect 6600 -1825 9305 -1775
use cc_inv  cc_inv_0
timestamp 1725397606
transform 1 0 65 0 1 40
box -60 -90 2805 1175
use cc_inv  cc_inv_1
timestamp 1725397606
transform 1 0 2930 0 1 40
box -60 -90 2805 1175
use cc_inv  cc_inv_2
timestamp 1725397606
transform 1 0 5795 0 1 40
box -60 -90 2805 1175
use cc_inv  cc_inv_3
timestamp 1725397606
transform -1 0 4615 0 -1 -650
box -60 -90 2805 1175
use cc_inv  cc_inv_4
timestamp 1725397606
transform -1 0 7480 0 -1 -650
box -60 -90 2805 1175
<< labels >>
rlabel metal1 1770 -1415 1770 -1415 1 OUT_P_0
port 3 n
rlabel metal1 1740 -890 1740 -890 1 OUT_n_0
port 4 n
rlabel space 2870 855 2870 855 1 OUT_P_1
port 5 n
rlabel space 2870 330 2870 330 1 OUT_N_1
port 6 n
rlabel space 5735 855 5735 855 1 OUT_P_2
port 7 n
rlabel space 5735 330 5735 330 1 OUT_N_2
port 8 n
rlabel metal1 8635 855 8635 855 1 OUT_P_3
port 9 n
rlabel metal1 8625 330 8625 330 1 OUT_N_3
port 10 n
rlabel space 4675 -890 4675 -890 1 OUT_N_4
port 11 n
rlabel space 4675 -1415 4675 -1415 1 OUT_P_4
port 12 n
<< end >>
