* NGSPICE file created from test_cc_inv.ext - technology: sky130A

.subckt test_main_inv A VPWR VGND Y VCCA GND
X0 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt test_aux_inv A VPWR VGND Y VCCA GND
X0 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt test_cc_inv IN_P IN_N VPWR VGND OUT_P OUT_N VCCA GND
Xtest_main_inv_0 IN_P VPWR VGND OUT_P VCCA GND test_main_inv
Xtest_main_inv_1 IN_N VPWR VGND OUT_N VCCA GND test_main_inv
Xtest_aux_inv_0 OUT_P VPWR VGND OUT_N VCCA GND test_aux_inv
Xtest_aux_inv_1 OUT_N VPWR VGND OUT_P VCCA GND test_aux_inv
.ends

