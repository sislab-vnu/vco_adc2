magic
tech sky130A
magscale 1 2
timestamp 1726742472
<< nwell >>
rect -808 1922 -430 1924
rect -832 1916 -522 1922
rect -832 1834 -564 1916
rect -832 1802 -546 1834
rect -832 1722 -570 1802
rect -812 1704 -570 1722
rect -566 1704 -546 1802
rect -812 1602 -258 1704
rect 972 1688 1024 1922
rect -840 1600 -258 1602
rect -1688 950 -1514 956
rect -1688 930 -1562 950
rect -1688 712 -1548 930
rect -1004 892 -800 956
rect -1004 872 -794 892
rect -656 872 -616 912
rect -1004 774 -994 872
rect -980 868 -794 872
rect -990 774 -794 868
rect -656 800 -616 840
rect -1004 760 -794 774
rect -1688 634 -1562 712
rect -1004 634 -800 760
rect -1688 632 -1476 634
<< pwell >>
rect -788 1496 -648 1502
rect -832 1360 -524 1496
rect 924 1360 1062 1428
rect -1014 1012 -760 1196
<< pdiff >>
rect -656 872 -616 912
rect -656 800 -616 840
<< psubdiff >>
rect -734 1428 -610 1442
rect -734 1394 -688 1428
rect -654 1394 -610 1428
rect -734 1380 -610 1394
rect -960 1112 -836 1126
rect -960 1078 -918 1112
rect -884 1078 -836 1112
rect -960 1064 -836 1078
<< nsubdiff >>
rect -632 1766 -570 1798
rect -632 1732 -618 1766
rect -584 1732 -570 1766
rect -632 1700 -570 1732
rect -1618 818 -1556 850
rect -1618 784 -1604 818
rect -1570 784 -1556 818
rect -1618 752 -1556 784
<< psubdiffcont >>
rect -688 1394 -654 1428
rect -918 1078 -884 1112
<< nsubdiffcont >>
rect -618 1732 -584 1766
rect -1604 784 -1570 818
<< locali >>
rect -632 1766 -570 1798
rect -632 1732 -618 1766
rect -584 1732 -570 1766
rect -632 1700 -570 1732
rect 856 1470 892 1504
rect -734 1428 -610 1442
rect -734 1394 -688 1428
rect -654 1394 -610 1428
rect 856 1402 892 1436
rect -734 1380 -610 1394
rect -960 1112 -836 1126
rect -960 1078 -918 1112
rect -884 1078 -836 1112
rect -960 1064 -836 1078
rect 840 1040 874 1062
rect 838 1034 880 1040
rect -1036 954 -651 1000
rect 838 998 840 1034
rect 874 998 880 1034
rect 838 970 880 998
rect -656 908 -616 912
rect -656 874 -654 908
rect -620 874 -616 908
rect -656 872 -616 874
rect -1618 818 -1556 850
rect -1618 784 -1604 818
rect -1570 784 -1556 818
rect -656 836 -616 840
rect -656 802 -654 836
rect -620 802 -616 836
rect -656 800 -616 802
rect -1618 752 -1556 784
<< viali >>
rect -618 1732 -584 1766
rect -1240 1552 -1200 1592
rect -882 1556 -848 1590
rect -508 1552 -468 1592
rect -250 1528 -216 1562
rect 856 1436 890 1470
rect -1380 972 -1346 1006
rect 840 998 874 1034
rect 1088 964 1132 1004
<< metal1 >>
rect -1438 2032 1480 2092
rect -1438 1604 -1390 2032
rect -632 1766 -570 1798
rect -632 1732 -618 1766
rect -584 1732 -570 1766
rect -632 1700 -570 1732
rect -1438 1592 -928 1604
rect -1438 1556 -1240 1592
rect -1252 1552 -1240 1556
rect -1200 1552 -928 1592
rect -1252 1540 -928 1552
rect -896 1600 -840 1676
rect -520 1600 -448 1664
rect -896 1592 -448 1600
rect -896 1590 -508 1592
rect -896 1556 -882 1590
rect -848 1556 -508 1590
rect -896 1552 -508 1556
rect -468 1552 -448 1592
rect -896 1544 -448 1552
rect -264 1562 -208 1600
rect -896 1502 -840 1544
rect -264 1528 -250 1562
rect -216 1528 -208 1562
rect -264 1502 -208 1528
rect -1842 1472 -208 1502
rect -1842 1010 -1802 1472
rect 840 1470 1320 1504
rect -734 1380 -610 1442
rect 840 1436 856 1470
rect 890 1444 1320 1470
rect 890 1436 908 1444
rect 840 1416 908 1436
rect -960 1064 -836 1126
rect 1260 1124 1320 1444
rect 828 1064 1320 1124
rect 828 1034 884 1064
rect -1410 1010 -1308 1012
rect -1842 1006 -1308 1010
rect -1842 972 -1380 1006
rect -1346 972 -1308 1006
rect -1842 970 -1308 972
rect -1410 952 -1308 970
rect 828 998 840 1034
rect 874 998 884 1034
rect 1420 1020 1480 2032
rect 828 958 884 998
rect 1072 1004 1480 1020
rect 1072 964 1088 1004
rect 1132 964 1480 1004
rect 1072 956 1480 964
rect 1072 892 1140 956
rect -1618 752 -1556 850
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform -1 0 -1004 0 -1 1216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_2  sky130_fd_sc_hd__dfxbp_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform -1 0 1158 0 -1 1216
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -538 0 1 1340
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -1274 0 1 1340
box -38 -48 498 592
<< end >>
