magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -260 -80 1660 1080
<< pwell >>
rect -106 -894 1646 -184
rect -246 -1036 1646 -894
rect -246 -1046 -114 -1036
<< nmos >>
rect 0 -1010 730 -210
rect 810 -1010 1540 -210
<< pmos >>
rect 0 0 730 1000
rect 810 0 1540 1000
<< ndiff >>
rect -80 -233 0 -210
rect -80 -267 -57 -233
rect -23 -267 0 -233
rect -80 -313 0 -267
rect -80 -347 -57 -313
rect -23 -347 0 -313
rect -80 -393 0 -347
rect -80 -427 -57 -393
rect -23 -427 0 -393
rect -80 -473 0 -427
rect -80 -507 -57 -473
rect -23 -507 0 -473
rect -80 -553 0 -507
rect -80 -587 -57 -553
rect -23 -587 0 -553
rect -80 -633 0 -587
rect -80 -667 -57 -633
rect -23 -667 0 -633
rect -80 -713 0 -667
rect -80 -747 -57 -713
rect -23 -747 0 -713
rect -80 -793 0 -747
rect -80 -827 -57 -793
rect -23 -827 0 -793
rect -80 -873 0 -827
rect -80 -907 -57 -873
rect -23 -907 0 -873
rect -80 -953 0 -907
rect -80 -987 -57 -953
rect -23 -987 0 -953
rect -80 -1010 0 -987
rect 730 -233 810 -210
rect 730 -267 753 -233
rect 787 -267 810 -233
rect 730 -313 810 -267
rect 730 -347 753 -313
rect 787 -347 810 -313
rect 730 -393 810 -347
rect 730 -427 753 -393
rect 787 -427 810 -393
rect 730 -473 810 -427
rect 730 -507 753 -473
rect 787 -507 810 -473
rect 730 -553 810 -507
rect 730 -587 753 -553
rect 787 -587 810 -553
rect 730 -633 810 -587
rect 730 -667 753 -633
rect 787 -667 810 -633
rect 730 -713 810 -667
rect 730 -747 753 -713
rect 787 -747 810 -713
rect 730 -793 810 -747
rect 730 -827 753 -793
rect 787 -827 810 -793
rect 730 -873 810 -827
rect 730 -907 753 -873
rect 787 -907 810 -873
rect 730 -953 810 -907
rect 730 -987 753 -953
rect 787 -987 810 -953
rect 730 -1010 810 -987
rect 1540 -233 1620 -210
rect 1540 -267 1563 -233
rect 1597 -267 1620 -233
rect 1540 -313 1620 -267
rect 1540 -347 1563 -313
rect 1597 -347 1620 -313
rect 1540 -393 1620 -347
rect 1540 -427 1563 -393
rect 1597 -427 1620 -393
rect 1540 -473 1620 -427
rect 1540 -507 1563 -473
rect 1597 -507 1620 -473
rect 1540 -553 1620 -507
rect 1540 -587 1563 -553
rect 1597 -587 1620 -553
rect 1540 -633 1620 -587
rect 1540 -667 1563 -633
rect 1597 -667 1620 -633
rect 1540 -713 1620 -667
rect 1540 -747 1563 -713
rect 1597 -747 1620 -713
rect 1540 -793 1620 -747
rect 1540 -827 1563 -793
rect 1597 -827 1620 -793
rect 1540 -873 1620 -827
rect 1540 -907 1563 -873
rect 1597 -907 1620 -873
rect 1540 -953 1620 -907
rect 1540 -987 1563 -953
rect 1597 -987 1620 -953
rect 1540 -1010 1620 -987
<< pdiff >>
rect -80 977 0 1000
rect -80 943 -57 977
rect -23 943 0 977
rect -80 897 0 943
rect -80 863 -57 897
rect -23 863 0 897
rect -80 817 0 863
rect -80 783 -57 817
rect -23 783 0 817
rect -80 737 0 783
rect -80 703 -57 737
rect -23 703 0 737
rect -80 657 0 703
rect -80 623 -57 657
rect -23 623 0 657
rect -80 577 0 623
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 730 977 810 1000
rect 730 943 753 977
rect 787 943 810 977
rect 730 897 810 943
rect 730 863 753 897
rect 787 863 810 897
rect 730 817 810 863
rect 730 783 753 817
rect 787 783 810 817
rect 730 737 810 783
rect 730 703 753 737
rect 787 703 810 737
rect 730 657 810 703
rect 730 623 753 657
rect 787 623 810 657
rect 730 577 810 623
rect 730 543 753 577
rect 787 543 810 577
rect 730 497 810 543
rect 730 463 753 497
rect 787 463 810 497
rect 730 417 810 463
rect 730 383 753 417
rect 787 383 810 417
rect 730 337 810 383
rect 730 303 753 337
rect 787 303 810 337
rect 730 257 810 303
rect 730 223 753 257
rect 787 223 810 257
rect 730 177 810 223
rect 730 143 753 177
rect 787 143 810 177
rect 730 97 810 143
rect 730 63 753 97
rect 787 63 810 97
rect 730 0 810 63
rect 1540 977 1620 1000
rect 1540 943 1563 977
rect 1597 943 1620 977
rect 1540 897 1620 943
rect 1540 863 1563 897
rect 1597 863 1620 897
rect 1540 817 1620 863
rect 1540 783 1563 817
rect 1597 783 1620 817
rect 1540 737 1620 783
rect 1540 703 1563 737
rect 1597 703 1620 737
rect 1540 657 1620 703
rect 1540 623 1563 657
rect 1597 623 1620 657
rect 1540 577 1620 623
rect 1540 543 1563 577
rect 1597 543 1620 577
rect 1540 497 1620 543
rect 1540 463 1563 497
rect 1597 463 1620 497
rect 1540 417 1620 463
rect 1540 383 1563 417
rect 1597 383 1620 417
rect 1540 337 1620 383
rect 1540 303 1563 337
rect 1597 303 1620 337
rect 1540 257 1620 303
rect 1540 223 1563 257
rect 1597 223 1620 257
rect 1540 177 1620 223
rect 1540 143 1563 177
rect 1597 143 1620 177
rect 1540 97 1620 143
rect 1540 63 1563 97
rect 1597 63 1620 97
rect 1540 0 1620 63
<< ndiffc >>
rect -57 -267 -23 -233
rect -57 -347 -23 -313
rect -57 -427 -23 -393
rect -57 -507 -23 -473
rect -57 -587 -23 -553
rect -57 -667 -23 -633
rect -57 -747 -23 -713
rect -57 -827 -23 -793
rect -57 -907 -23 -873
rect -57 -987 -23 -953
rect 753 -267 787 -233
rect 753 -347 787 -313
rect 753 -427 787 -393
rect 753 -507 787 -473
rect 753 -587 787 -553
rect 753 -667 787 -633
rect 753 -747 787 -713
rect 753 -827 787 -793
rect 753 -907 787 -873
rect 753 -987 787 -953
rect 1563 -267 1597 -233
rect 1563 -347 1597 -313
rect 1563 -427 1597 -393
rect 1563 -507 1597 -473
rect 1563 -587 1597 -553
rect 1563 -667 1597 -633
rect 1563 -747 1597 -713
rect 1563 -827 1597 -793
rect 1563 -907 1597 -873
rect 1563 -987 1597 -953
<< pdiffc >>
rect -57 943 -23 977
rect -57 863 -23 897
rect -57 783 -23 817
rect -57 703 -23 737
rect -57 623 -23 657
rect -57 543 -23 577
rect -57 463 -23 497
rect -57 383 -23 417
rect -57 303 -23 337
rect -57 223 -23 257
rect -57 143 -23 177
rect -57 63 -23 97
rect 753 943 787 977
rect 753 863 787 897
rect 753 783 787 817
rect 753 703 787 737
rect 753 623 787 657
rect 753 543 787 577
rect 753 463 787 497
rect 753 383 787 417
rect 753 303 787 337
rect 753 223 787 257
rect 753 143 787 177
rect 753 63 787 97
rect 1563 943 1597 977
rect 1563 863 1597 897
rect 1563 783 1597 817
rect 1563 703 1597 737
rect 1563 623 1597 657
rect 1563 543 1597 577
rect 1563 463 1597 497
rect 1563 383 1597 417
rect 1563 303 1597 337
rect 1563 223 1597 257
rect 1563 143 1597 177
rect 1563 63 1597 97
<< psubdiff >>
rect -220 -953 -140 -920
rect -220 -987 -197 -953
rect -163 -987 -140 -953
rect -220 -1020 -140 -987
<< nsubdiff >>
rect -220 977 -140 1010
rect -220 943 -197 977
rect -163 943 -140 977
rect -220 910 -140 943
<< psubdiffcont >>
rect -197 -987 -163 -953
<< nsubdiffcont >>
rect -197 943 -163 977
<< poly >>
rect 0 1000 730 1080
rect 810 1000 1540 1080
rect 0 -30 730 0
rect 810 -30 1540 0
rect 0 -93 1540 -30
rect 0 -127 183 -93
rect 217 -127 263 -93
rect 297 -127 343 -93
rect 377 -127 923 -93
rect 957 -127 1003 -93
rect 1037 -127 1083 -93
rect 1117 -127 1540 -93
rect 0 -180 1540 -127
rect 0 -210 730 -180
rect 810 -210 1540 -180
rect 0 -1090 730 -1010
rect 810 -1090 1540 -1010
<< polycont >>
rect 183 -127 217 -93
rect 263 -127 297 -93
rect 343 -127 377 -93
rect 923 -127 957 -93
rect 1003 -127 1037 -93
rect 1083 -127 1117 -93
<< locali >>
rect -80 1180 1620 1260
rect -220 977 -140 1010
rect -220 943 -197 977
rect -163 943 -140 977
rect -220 910 -140 943
rect -80 977 0 1180
rect -80 943 -57 977
rect -23 943 0 977
rect -80 897 0 943
rect -80 863 -57 897
rect -23 863 0 897
rect -80 817 0 863
rect -80 783 -57 817
rect -23 783 0 817
rect -80 737 0 783
rect -80 703 -57 737
rect -23 703 0 737
rect -80 657 0 703
rect -80 623 -57 657
rect -23 623 0 657
rect -80 577 0 623
rect -80 543 -57 577
rect -23 543 0 577
rect -80 497 0 543
rect -80 463 -57 497
rect -23 463 0 497
rect -80 417 0 463
rect -80 383 -57 417
rect -23 383 0 417
rect -80 337 0 383
rect -80 303 -57 337
rect -23 303 0 337
rect -80 257 0 303
rect -80 223 -57 257
rect -23 223 0 257
rect -80 177 0 223
rect -80 143 -57 177
rect -23 143 0 177
rect -80 97 0 143
rect -80 63 -57 97
rect -23 63 0 97
rect -80 0 0 63
rect 730 977 810 1000
rect 730 943 753 977
rect 787 943 810 977
rect 730 897 810 943
rect 730 863 753 897
rect 787 863 810 897
rect 730 817 810 863
rect 730 783 753 817
rect 787 783 810 817
rect 730 737 810 783
rect 730 703 753 737
rect 787 703 810 737
rect 730 657 810 703
rect 730 623 753 657
rect 787 623 810 657
rect 730 577 810 623
rect 730 543 753 577
rect 787 543 810 577
rect 730 497 810 543
rect 730 463 753 497
rect 787 463 810 497
rect 730 417 810 463
rect 730 383 753 417
rect 787 383 810 417
rect 730 337 810 383
rect 730 303 753 337
rect 787 303 810 337
rect 730 257 810 303
rect 730 223 753 257
rect 787 223 810 257
rect 730 177 810 223
rect 730 143 753 177
rect 787 143 810 177
rect 730 97 810 143
rect 730 63 753 97
rect 787 63 810 97
rect 160 -93 400 -40
rect 160 -127 183 -93
rect 217 -127 263 -93
rect 297 -127 343 -93
rect 377 -127 400 -93
rect 160 -170 400 -127
rect -80 -233 0 -210
rect -80 -267 -57 -233
rect -23 -267 0 -233
rect -80 -313 0 -267
rect -80 -347 -57 -313
rect -23 -347 0 -313
rect -80 -393 0 -347
rect -80 -427 -57 -393
rect -23 -427 0 -393
rect -80 -473 0 -427
rect -80 -507 -57 -473
rect -23 -507 0 -473
rect -80 -553 0 -507
rect -80 -587 -57 -553
rect -23 -587 0 -553
rect -80 -633 0 -587
rect -80 -667 -57 -633
rect -23 -667 0 -633
rect -80 -713 0 -667
rect -80 -747 -57 -713
rect -23 -747 0 -713
rect -80 -793 0 -747
rect -80 -827 -57 -793
rect -23 -827 0 -793
rect -80 -873 0 -827
rect -80 -907 -57 -873
rect -23 -907 0 -873
rect -220 -953 -140 -920
rect -220 -987 -197 -953
rect -163 -987 -140 -953
rect -220 -1020 -140 -987
rect -80 -953 0 -907
rect -80 -987 -57 -953
rect -23 -987 0 -953
rect -80 -1190 0 -987
rect 730 -233 810 63
rect 1540 977 1620 1180
rect 1540 943 1563 977
rect 1597 943 1620 977
rect 1540 897 1620 943
rect 1540 863 1563 897
rect 1597 863 1620 897
rect 1540 817 1620 863
rect 1540 783 1563 817
rect 1597 783 1620 817
rect 1540 737 1620 783
rect 1540 703 1563 737
rect 1597 703 1620 737
rect 1540 657 1620 703
rect 1540 623 1563 657
rect 1597 623 1620 657
rect 1540 577 1620 623
rect 1540 543 1563 577
rect 1597 543 1620 577
rect 1540 497 1620 543
rect 1540 463 1563 497
rect 1597 463 1620 497
rect 1540 417 1620 463
rect 1540 383 1563 417
rect 1597 383 1620 417
rect 1540 337 1620 383
rect 1540 303 1563 337
rect 1597 303 1620 337
rect 1540 257 1620 303
rect 1540 223 1563 257
rect 1597 223 1620 257
rect 1540 177 1620 223
rect 1540 143 1563 177
rect 1597 143 1620 177
rect 1540 97 1620 143
rect 1540 63 1563 97
rect 1597 63 1620 97
rect 1540 0 1620 63
rect 900 -93 1140 -40
rect 900 -127 923 -93
rect 957 -127 1003 -93
rect 1037 -127 1083 -93
rect 1117 -127 1140 -93
rect 900 -170 1140 -127
rect 730 -267 753 -233
rect 787 -267 810 -233
rect 730 -313 810 -267
rect 730 -347 753 -313
rect 787 -347 810 -313
rect 730 -393 810 -347
rect 730 -427 753 -393
rect 787 -427 810 -393
rect 730 -473 810 -427
rect 730 -507 753 -473
rect 787 -507 810 -473
rect 730 -553 810 -507
rect 730 -587 753 -553
rect 787 -587 810 -553
rect 730 -633 810 -587
rect 730 -667 753 -633
rect 787 -667 810 -633
rect 730 -713 810 -667
rect 730 -747 753 -713
rect 787 -747 810 -713
rect 730 -793 810 -747
rect 730 -827 753 -793
rect 787 -827 810 -793
rect 730 -873 810 -827
rect 730 -907 753 -873
rect 787 -907 810 -873
rect 730 -953 810 -907
rect 730 -987 753 -953
rect 787 -987 810 -953
rect 730 -1010 810 -987
rect 1540 -233 1620 -210
rect 1540 -267 1563 -233
rect 1597 -267 1620 -233
rect 1540 -313 1620 -267
rect 1540 -347 1563 -313
rect 1597 -347 1620 -313
rect 1540 -393 1620 -347
rect 1540 -427 1563 -393
rect 1597 -427 1620 -393
rect 1540 -473 1620 -427
rect 1540 -507 1563 -473
rect 1597 -507 1620 -473
rect 1540 -553 1620 -507
rect 1540 -587 1563 -553
rect 1597 -587 1620 -553
rect 1540 -633 1620 -587
rect 1540 -667 1563 -633
rect 1597 -667 1620 -633
rect 1540 -713 1620 -667
rect 1540 -747 1563 -713
rect 1597 -747 1620 -713
rect 1540 -793 1620 -747
rect 1540 -827 1563 -793
rect 1597 -827 1620 -793
rect 1540 -873 1620 -827
rect 1540 -907 1563 -873
rect 1597 -907 1620 -873
rect 1540 -953 1620 -907
rect 1540 -987 1563 -953
rect 1597 -987 1620 -953
rect 1540 -1190 1620 -987
rect -80 -1270 1620 -1190
<< viali >>
rect -197 943 -163 977
rect 183 -127 217 -93
rect 263 -127 297 -93
rect 343 -127 377 -93
rect -197 -987 -163 -953
rect 923 -127 957 -93
rect 1003 -127 1037 -93
rect 1083 -127 1117 -93
<< metal1 >>
rect -220 977 -140 1010
rect -220 943 -197 977
rect -163 943 -140 977
rect -220 910 -140 943
rect 160 -93 1140 -40
rect 160 -127 183 -93
rect 217 -127 263 -93
rect 297 -127 343 -93
rect 377 -127 923 -93
rect 957 -127 1003 -93
rect 1037 -127 1083 -93
rect 1117 -127 1140 -93
rect 160 -170 1140 -127
rect -220 -953 -140 -920
rect -220 -987 -197 -953
rect -163 -987 -140 -953
rect -220 -1020 -140 -987
<< labels >>
rlabel metal1 s 160 -110 160 -110 4 A
rlabel locali s 770 1260 770 1260 4 VPWR
rlabel locali s 770 -1270 770 -1270 4 VGND
rlabel locali s 770 -1010 770 -1010 4 Y
rlabel metal1 s -180 1010 -180 1010 4 VCCA
rlabel metal1 s -180 -1020 -180 -1020 4 GND
<< end >>
