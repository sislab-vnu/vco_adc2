magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< poly >>
rect -48 614 48 630
rect -48 580 -17 614
rect 17 580 48 614
rect -48 200 48 580
rect -48 -580 48 -200
rect -48 -614 -17 -580
rect 17 -614 48 -580
rect -48 -630 48 -614
<< polycont >>
rect -17 580 17 614
rect -17 -614 17 -580
<< npolyres >>
rect -48 -200 48 200
<< locali >>
rect -48 580 -17 614
rect 17 580 48 614
rect -32 578 -17 580
rect 17 578 32 580
rect -32 540 32 578
rect -32 506 -17 540
rect 17 506 32 540
rect -32 468 32 506
rect -32 434 -17 468
rect 17 434 32 468
rect -32 396 32 434
rect -32 362 -17 396
rect 17 362 32 396
rect -32 324 32 362
rect -32 290 -17 324
rect 17 290 32 324
rect -32 252 32 290
rect -32 218 -17 252
rect 17 218 32 252
rect -32 217 32 218
rect -32 -219 32 -217
rect -32 -253 -17 -219
rect 17 -253 32 -219
rect -32 -291 32 -253
rect -32 -325 -17 -291
rect 17 -325 32 -291
rect -32 -363 32 -325
rect -32 -397 -17 -363
rect 17 -397 32 -363
rect -32 -435 32 -397
rect -32 -469 -17 -435
rect 17 -469 32 -435
rect -32 -507 32 -469
rect -32 -541 -17 -507
rect 17 -541 32 -507
rect -32 -579 32 -541
rect -32 -580 -17 -579
rect 17 -580 32 -579
rect -48 -614 -17 -580
rect 17 -614 48 -580
<< viali >>
rect -17 580 17 612
rect -17 578 17 580
rect -17 506 17 540
rect -17 434 17 468
rect -17 362 17 396
rect -17 290 17 324
rect -17 218 17 252
rect -17 -253 17 -219
rect -17 -325 17 -291
rect -17 -397 17 -363
rect -17 -469 17 -435
rect -17 -541 17 -507
rect -17 -580 17 -579
rect -17 -613 17 -580
<< metal1 >>
rect -38 612 38 626
rect -38 578 -17 612
rect 17 578 38 612
rect -38 540 38 578
rect -38 506 -17 540
rect 17 506 38 540
rect -38 468 38 506
rect -38 434 -17 468
rect 17 434 38 468
rect -38 396 38 434
rect -38 362 -17 396
rect 17 362 38 396
rect -38 324 38 362
rect -38 290 -17 324
rect 17 290 38 324
rect -38 252 38 290
rect -38 218 -17 252
rect 17 218 38 252
rect -38 205 38 218
rect -38 -219 38 -205
rect -38 -253 -17 -219
rect 17 -253 38 -219
rect -38 -291 38 -253
rect -38 -325 -17 -291
rect 17 -325 38 -291
rect -38 -363 38 -325
rect -38 -397 -17 -363
rect 17 -397 38 -363
rect -38 -435 38 -397
rect -38 -469 -17 -435
rect 17 -469 38 -435
rect -38 -507 38 -469
rect -38 -541 -17 -507
rect 17 -541 38 -507
rect -38 -579 38 -541
rect -38 -613 -17 -579
rect 17 -613 38 -579
rect -38 -626 38 -613
<< end >>
