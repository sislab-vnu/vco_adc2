VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 109.180 3381.220 112.680 3381.320 ;
        RECT 107.365 3380.900 112.680 3381.220 ;
        RECT 109.180 3380.620 112.680 3380.900 ;
      LAYER met1 ;
        RECT 112.630 3381.320 113.880 3381.420 ;
        RECT 107.305 3380.870 109.410 3381.250 ;
        RECT 111.680 3380.620 113.880 3381.320 ;
      LAYER met2 ;
        RECT 283.770 3518.770 284.330 3524.800 ;
        RECT 275.750 3516.930 286.330 3518.770 ;
        RECT 275.630 3382.120 277.630 3516.930 ;
        RECT 181.180 3381.620 277.630 3382.120 ;
        RECT 113.880 3381.420 277.630 3381.620 ;
        RECT 112.630 3380.620 277.630 3381.420 ;
        RECT 181.180 3380.120 277.630 3380.620 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 117.080 3330.970 117.380 3331.470 ;
        RECT 131.630 3330.920 132.130 3331.420 ;
      LAYER met1 ;
        RECT 113.180 3334.120 114.280 3334.620 ;
        RECT 113.180 3333.620 132.130 3334.120 ;
        RECT 113.180 3333.520 114.280 3333.620 ;
        RECT 118.430 3331.470 118.930 3333.620 ;
        RECT 116.880 3330.970 118.930 3331.470 ;
        RECT 131.630 3330.920 132.130 3333.620 ;
      LAYER met2 ;
        RECT 1.000 3486.970 9.160 3488.880 ;
        RECT 1.000 3484.970 44.030 3486.970 ;
        RECT 1.000 3484.120 9.160 3484.970 ;
        RECT 42.030 3369.570 44.030 3484.970 ;
        RECT 42.030 3368.470 93.680 3369.570 ;
        RECT 92.580 3358.420 93.680 3368.470 ;
        RECT 92.580 3357.320 103.280 3358.420 ;
        RECT 102.180 3334.620 103.280 3357.320 ;
        RECT 102.180 3333.520 114.280 3334.620 ;
      LAYER met3 ;
        RECT 1.000 3487.300 9.160 3488.880 ;
        RECT -4.800 3486.100 9.160 3487.300 ;
        RECT 1.000 3484.120 9.160 3486.100 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER li1 ;
        RECT 120.830 3330.970 121.830 3331.470 ;
        RECT 126.130 3330.970 128.430 3331.470 ;
      LAYER met1 ;
        RECT 123.730 3331.470 124.730 3331.970 ;
        RECT 120.630 3330.970 128.430 3331.470 ;
      LAYER met2 ;
        RECT 16.080 3337.620 100.880 3338.620 ;
        RECT 1.000 3225.770 9.160 3227.760 ;
        RECT 16.080 3225.770 18.080 3337.620 ;
        RECT 99.880 3326.370 100.880 3337.620 ;
        RECT 123.730 3328.020 124.730 3331.970 ;
        RECT 114.180 3327.020 124.730 3328.020 ;
        RECT 114.180 3326.370 115.180 3327.020 ;
        RECT 99.880 3325.370 115.180 3326.370 ;
        RECT 1.000 3223.770 18.080 3225.770 ;
        RECT 1.000 3223.000 9.160 3223.770 ;
      LAYER met3 ;
        RECT 1.000 3226.180 9.160 3227.760 ;
        RECT -4.800 3224.980 9.160 3226.180 ;
        RECT 1.000 3223.000 9.160 3224.980 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 65.770 2873.810 65.780 ;
        RECT 2859.820 65.470 2873.810 65.770 ;
        RECT 2873.430 65.460 2873.810 65.470 ;
        RECT 2873.430 33.130 2873.810 33.140 ;
        RECT 2917.600 33.130 2924.800 33.580 ;
        RECT 2873.430 32.830 2924.800 33.130 ;
        RECT 2873.430 32.820 2873.810 32.830 ;
        RECT 2917.600 32.380 2924.800 32.830 ;
      LAYER met4 ;
        RECT 2873.455 65.455 2873.785 65.785 ;
        RECT 2873.470 33.145 2873.770 65.455 ;
        RECT 2873.455 32.815 2873.785 33.145 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 282.010 2873.810 282.020 ;
        RECT 2859.820 281.710 2873.810 282.010 ;
        RECT 2873.430 281.700 2873.810 281.710 ;
        RECT 2873.430 231.690 2873.810 231.700 ;
        RECT 2917.600 231.690 2924.800 232.140 ;
        RECT 2873.430 231.390 2924.800 231.690 ;
        RECT 2873.430 231.380 2873.810 231.390 ;
        RECT 2917.600 230.940 2924.800 231.390 ;
      LAYER met4 ;
        RECT 2873.455 281.695 2873.785 282.025 ;
        RECT 2873.470 231.705 2873.770 281.695 ;
        RECT 2873.455 231.375 2873.785 231.705 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 498.250 2874.730 498.260 ;
        RECT 2859.820 497.950 2874.730 498.250 ;
        RECT 2874.350 497.940 2874.730 497.950 ;
        RECT 2874.350 430.930 2874.730 430.940 ;
        RECT 2917.600 430.930 2924.800 431.380 ;
        RECT 2874.350 430.630 2924.800 430.930 ;
        RECT 2874.350 430.620 2874.730 430.630 ;
        RECT 2917.600 430.180 2924.800 430.630 ;
      LAYER met4 ;
        RECT 2874.375 497.935 2874.705 498.265 ;
        RECT 2874.390 430.945 2874.690 497.935 ;
        RECT 2874.375 430.615 2874.705 430.945 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.890 2.400 1857.340 ;
        RECT 18.670 1856.890 19.050 1856.900 ;
        RECT -4.800 1856.590 19.050 1856.890 ;
        RECT -4.800 1856.140 2.400 1856.590 ;
        RECT 18.670 1856.580 19.050 1856.590 ;
        RECT 18.670 1723.610 19.050 1723.620 ;
        RECT 18.670 1723.310 60.260 1723.610 ;
        RECT 18.670 1723.300 19.050 1723.310 ;
      LAYER met4 ;
        RECT 18.695 1856.575 19.025 1856.905 ;
        RECT 18.710 1723.625 19.010 1856.575 ;
        RECT 18.695 1723.295 19.025 1723.625 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1596.450 2.400 1596.900 ;
        RECT 18.670 1596.450 19.050 1596.460 ;
        RECT -4.800 1596.150 19.050 1596.450 ;
        RECT -4.800 1595.700 2.400 1596.150 ;
        RECT 18.670 1596.140 19.050 1596.150 ;
        RECT 18.670 1507.370 19.050 1507.380 ;
        RECT 18.670 1507.070 60.260 1507.370 ;
        RECT 18.670 1507.060 19.050 1507.070 ;
      LAYER met4 ;
        RECT 18.695 1596.135 19.025 1596.465 ;
        RECT 18.710 1507.385 19.010 1596.135 ;
        RECT 18.695 1507.055 19.025 1507.385 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1336.010 2.400 1336.460 ;
        RECT 40.750 1336.010 41.130 1336.020 ;
        RECT -4.800 1335.710 41.130 1336.010 ;
        RECT -4.800 1335.260 2.400 1335.710 ;
        RECT 40.750 1335.700 41.130 1335.710 ;
        RECT 40.750 1291.130 41.130 1291.140 ;
        RECT 40.750 1290.830 60.260 1291.130 ;
        RECT 40.750 1290.820 41.130 1290.830 ;
      LAYER met4 ;
        RECT 40.775 1335.695 41.105 1336.025 ;
        RECT 40.790 1291.145 41.090 1335.695 ;
        RECT 40.775 1290.815 41.105 1291.145 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.890 2.400 1075.340 ;
        RECT -4.800 1074.590 60.260 1074.890 ;
        RECT -4.800 1074.140 2.400 1074.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.550 858.650 31.930 858.660 ;
        RECT 31.550 858.350 60.260 858.650 ;
        RECT 31.550 858.340 31.930 858.350 ;
        RECT -4.800 814.450 2.400 814.900 ;
        RECT 31.550 814.450 31.930 814.460 ;
        RECT -4.800 814.150 31.930 814.450 ;
        RECT -4.800 813.700 2.400 814.150 ;
        RECT 31.550 814.140 31.930 814.150 ;
      LAYER met4 ;
        RECT 31.575 858.335 31.905 858.665 ;
        RECT 31.590 814.465 31.890 858.335 ;
        RECT 31.575 814.135 31.905 814.465 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.830 642.410 17.210 642.420 ;
        RECT 16.830 642.110 60.260 642.410 ;
        RECT 16.830 642.100 17.210 642.110 ;
        RECT -4.800 553.330 2.400 553.780 ;
        RECT 16.830 553.330 17.210 553.340 ;
        RECT -4.800 553.030 17.210 553.330 ;
        RECT -4.800 552.580 2.400 553.030 ;
        RECT 16.830 553.020 17.210 553.030 ;
      LAYER met4 ;
        RECT 16.855 642.095 17.185 642.425 ;
        RECT 16.870 553.345 17.170 642.095 ;
        RECT 16.855 553.015 17.185 553.345 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 43.510 426.170 43.890 426.180 ;
        RECT 43.510 425.870 60.260 426.170 ;
        RECT 43.510 425.860 43.890 425.870 ;
        RECT -4.800 358.170 2.400 358.620 ;
        RECT 43.510 358.170 43.890 358.180 ;
        RECT -4.800 357.870 43.890 358.170 ;
        RECT -4.800 357.420 2.400 357.870 ;
        RECT 43.510 357.860 43.890 357.870 ;
      LAYER met4 ;
        RECT 43.535 425.855 43.865 426.185 ;
        RECT 43.550 358.185 43.850 425.855 ;
        RECT 43.535 357.855 43.865 358.185 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.430 209.930 44.810 209.940 ;
        RECT 44.430 209.630 60.260 209.930 ;
        RECT 44.430 209.620 44.810 209.630 ;
        RECT -4.800 162.330 2.400 162.780 ;
        RECT 44.430 162.330 44.810 162.340 ;
        RECT -4.800 162.030 44.810 162.330 ;
        RECT -4.800 161.580 2.400 162.030 ;
        RECT 44.430 162.020 44.810 162.030 ;
      LAYER met4 ;
        RECT 44.455 209.615 44.785 209.945 ;
        RECT 44.470 162.345 44.770 209.615 ;
        RECT 44.455 162.015 44.785 162.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 714.490 2873.810 714.500 ;
        RECT 2859.820 714.190 2873.810 714.490 ;
        RECT 2873.430 714.180 2873.810 714.190 ;
        RECT 2873.430 630.170 2873.810 630.180 ;
        RECT 2917.600 630.170 2924.800 630.620 ;
        RECT 2873.430 629.870 2924.800 630.170 ;
        RECT 2873.430 629.860 2873.810 629.870 ;
        RECT 2917.600 629.420 2924.800 629.870 ;
      LAYER met4 ;
        RECT 2873.455 714.175 2873.785 714.505 ;
        RECT 2873.470 630.185 2873.770 714.175 ;
        RECT 2873.455 629.855 2873.785 630.185 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 930.730 2874.730 930.740 ;
        RECT 2859.820 930.430 2874.730 930.730 ;
        RECT 2874.350 930.420 2874.730 930.430 ;
        RECT 2874.350 829.410 2874.730 829.420 ;
        RECT 2917.600 829.410 2924.800 829.860 ;
        RECT 2874.350 829.110 2924.800 829.410 ;
        RECT 2874.350 829.100 2874.730 829.110 ;
        RECT 2917.600 828.660 2924.800 829.110 ;
      LAYER met4 ;
        RECT 2874.375 930.415 2874.705 930.745 ;
        RECT 2874.390 829.425 2874.690 930.415 ;
        RECT 2874.375 829.095 2874.705 829.425 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 1146.970 2873.810 1146.980 ;
        RECT 2859.820 1146.670 2873.810 1146.970 ;
        RECT 2873.430 1146.660 2873.810 1146.670 ;
        RECT 2873.430 1028.650 2873.810 1028.660 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2873.430 1028.350 2924.800 1028.650 ;
        RECT 2873.430 1028.340 2873.810 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
      LAYER met4 ;
        RECT 2873.455 1146.655 2873.785 1146.985 ;
        RECT 2873.470 1028.665 2873.770 1146.655 ;
        RECT 2873.455 1028.335 2873.785 1028.665 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 1363.210 2874.730 1363.220 ;
        RECT 2859.820 1362.910 2874.730 1363.210 ;
        RECT 2874.350 1362.900 2874.730 1362.910 ;
        RECT 2874.350 1227.890 2874.730 1227.900 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2874.350 1227.590 2924.800 1227.890 ;
        RECT 2874.350 1227.580 2874.730 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
      LAYER met4 ;
        RECT 2874.375 1362.895 2874.705 1363.225 ;
        RECT 2874.390 1227.905 2874.690 1362.895 ;
        RECT 2874.375 1227.575 2874.705 1227.905 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2875.270 1579.450 2875.650 1579.460 ;
        RECT 2859.820 1579.150 2875.650 1579.450 ;
        RECT 2875.270 1579.140 2875.650 1579.150 ;
        RECT 2875.270 1493.770 2875.650 1493.780 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2875.270 1493.470 2924.800 1493.770 ;
        RECT 2875.270 1493.460 2875.650 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
      LAYER met4 ;
        RECT 2875.295 1579.135 2875.625 1579.465 ;
        RECT 2875.310 1493.785 2875.610 1579.135 ;
        RECT 2875.295 1493.455 2875.625 1493.785 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 209.930 2873.810 209.940 ;
        RECT 2859.820 209.630 2873.810 209.930 ;
        RECT 2873.430 209.620 2873.810 209.630 ;
        RECT 2873.430 165.730 2873.810 165.740 ;
        RECT 2917.600 165.730 2924.800 166.180 ;
        RECT 2873.430 165.430 2924.800 165.730 ;
        RECT 2873.430 165.420 2873.810 165.430 ;
        RECT 2917.600 164.980 2924.800 165.430 ;
      LAYER met4 ;
        RECT 2873.455 209.615 2873.785 209.945 ;
        RECT 2873.470 165.745 2873.770 209.615 ;
        RECT 2873.455 165.415 2873.785 165.745 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 426.170 2873.810 426.180 ;
        RECT 2859.820 425.870 2873.810 426.170 ;
        RECT 2873.430 425.860 2873.810 425.870 ;
        RECT 2873.430 364.970 2873.810 364.980 ;
        RECT 2917.600 364.970 2924.800 365.420 ;
        RECT 2873.430 364.670 2924.800 364.970 ;
        RECT 2873.430 364.660 2873.810 364.670 ;
        RECT 2917.600 364.220 2924.800 364.670 ;
      LAYER met4 ;
        RECT 2873.455 425.855 2873.785 426.185 ;
        RECT 2873.470 364.985 2873.770 425.855 ;
        RECT 2873.455 364.655 2873.785 364.985 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 642.410 2874.730 642.420 ;
        RECT 2859.820 642.110 2874.730 642.410 ;
        RECT 2874.350 642.100 2874.730 642.110 ;
        RECT 2874.350 564.210 2874.730 564.220 ;
        RECT 2917.600 564.210 2924.800 564.660 ;
        RECT 2874.350 563.910 2924.800 564.210 ;
        RECT 2874.350 563.900 2874.730 563.910 ;
        RECT 2917.600 563.460 2924.800 563.910 ;
      LAYER met4 ;
        RECT 2874.375 642.095 2874.705 642.425 ;
        RECT 2874.390 564.225 2874.690 642.095 ;
        RECT 2874.375 563.895 2874.705 564.225 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1727.010 2.400 1727.460 ;
        RECT 16.830 1727.010 17.210 1727.020 ;
        RECT -4.800 1726.710 17.210 1727.010 ;
        RECT -4.800 1726.260 2.400 1726.710 ;
        RECT 16.830 1726.700 17.210 1726.710 ;
        RECT 16.830 1579.450 17.210 1579.460 ;
        RECT 16.830 1579.150 60.260 1579.450 ;
        RECT 16.830 1579.140 17.210 1579.150 ;
      LAYER met4 ;
        RECT 16.855 1726.695 17.185 1727.025 ;
        RECT 16.870 1579.465 17.170 1726.695 ;
        RECT 16.855 1579.135 17.185 1579.465 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.890 2.400 1466.340 ;
        RECT 16.830 1465.890 17.210 1465.900 ;
        RECT -4.800 1465.590 17.210 1465.890 ;
        RECT -4.800 1465.140 2.400 1465.590 ;
        RECT 16.830 1465.580 17.210 1465.590 ;
        RECT 16.830 1363.210 17.210 1363.220 ;
        RECT 16.830 1362.910 60.260 1363.210 ;
        RECT 16.830 1362.900 17.210 1362.910 ;
      LAYER met4 ;
        RECT 16.855 1465.575 17.185 1465.905 ;
        RECT 16.870 1363.225 17.170 1465.575 ;
        RECT 16.855 1362.895 17.185 1363.225 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1205.450 2.400 1205.900 ;
        RECT 37.070 1205.450 37.450 1205.460 ;
        RECT -4.800 1205.150 37.450 1205.450 ;
        RECT -4.800 1204.700 2.400 1205.150 ;
        RECT 37.070 1205.140 37.450 1205.150 ;
        RECT 37.070 1146.970 37.450 1146.980 ;
        RECT 37.070 1146.670 60.260 1146.970 ;
        RECT 37.070 1146.660 37.450 1146.670 ;
      LAYER met4 ;
        RECT 37.095 1205.135 37.425 1205.465 ;
        RECT 37.110 1146.985 37.410 1205.135 ;
        RECT 37.095 1146.655 37.425 1146.985 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 944.330 2.400 944.780 ;
        RECT 31.550 944.330 31.930 944.340 ;
        RECT -4.800 944.030 31.930 944.330 ;
        RECT -4.800 943.580 2.400 944.030 ;
        RECT 31.550 944.020 31.930 944.030 ;
        RECT 31.550 930.730 31.930 930.740 ;
        RECT 31.550 930.430 60.260 930.730 ;
        RECT 31.550 930.420 31.930 930.430 ;
      LAYER met4 ;
        RECT 31.575 944.015 31.905 944.345 ;
        RECT 31.590 930.745 31.890 944.015 ;
        RECT 31.575 930.415 31.905 930.745 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.190 714.490 24.570 714.500 ;
        RECT 24.190 714.190 60.260 714.490 ;
        RECT 24.190 714.180 24.570 714.190 ;
        RECT -4.800 683.890 2.400 684.340 ;
        RECT 24.190 683.890 24.570 683.900 ;
        RECT -4.800 683.590 24.570 683.890 ;
        RECT -4.800 683.140 2.400 683.590 ;
        RECT 24.190 683.580 24.570 683.590 ;
      LAYER met4 ;
        RECT 24.215 714.175 24.545 714.505 ;
        RECT 24.230 683.905 24.530 714.175 ;
        RECT 24.215 683.575 24.545 683.905 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.430 498.250 44.810 498.260 ;
        RECT 44.430 497.950 60.260 498.250 ;
        RECT 44.430 497.940 44.810 497.950 ;
        RECT -4.800 423.450 2.400 423.900 ;
        RECT 44.430 423.450 44.810 423.460 ;
        RECT -4.800 423.150 44.810 423.450 ;
        RECT -4.800 422.700 2.400 423.150 ;
        RECT 44.430 423.140 44.810 423.150 ;
      LAYER met4 ;
        RECT 44.455 497.935 44.785 498.265 ;
        RECT 44.470 423.465 44.770 497.935 ;
        RECT 44.455 423.135 44.785 423.465 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.430 282.010 44.810 282.020 ;
        RECT 44.430 281.710 60.260 282.010 ;
        RECT 44.430 281.700 44.810 281.710 ;
        RECT -4.800 227.610 2.400 228.060 ;
        RECT 44.430 227.610 44.810 227.620 ;
        RECT -4.800 227.310 44.810 227.610 ;
        RECT -4.800 226.860 2.400 227.310 ;
        RECT 44.430 227.300 44.810 227.310 ;
      LAYER met4 ;
        RECT 44.455 281.695 44.785 282.025 ;
        RECT 44.470 227.625 44.770 281.695 ;
        RECT 44.455 227.295 44.785 227.625 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.430 65.770 44.810 65.780 ;
        RECT 44.430 65.470 60.260 65.770 ;
        RECT 44.430 65.460 44.810 65.470 ;
        RECT -4.800 32.450 2.400 32.900 ;
        RECT 44.430 32.450 44.810 32.460 ;
        RECT -4.800 32.150 44.810 32.450 ;
        RECT -4.800 31.700 2.400 32.150 ;
        RECT 44.430 32.140 44.810 32.150 ;
      LAYER met4 ;
        RECT 44.455 65.455 44.785 65.785 ;
        RECT 44.470 32.465 44.770 65.455 ;
        RECT 44.455 32.135 44.785 32.465 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 858.650 2873.810 858.660 ;
        RECT 2859.820 858.350 2873.810 858.650 ;
        RECT 2873.430 858.340 2873.810 858.350 ;
        RECT 2873.430 763.450 2873.810 763.460 ;
        RECT 2917.600 763.450 2924.800 763.900 ;
        RECT 2873.430 763.150 2924.800 763.450 ;
        RECT 2873.430 763.140 2873.810 763.150 ;
        RECT 2917.600 762.700 2924.800 763.150 ;
      LAYER met4 ;
        RECT 2873.455 858.335 2873.785 858.665 ;
        RECT 2873.470 763.465 2873.770 858.335 ;
        RECT 2873.455 763.135 2873.785 763.465 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 1074.890 2874.730 1074.900 ;
        RECT 2859.820 1074.590 2874.730 1074.890 ;
        RECT 2874.350 1074.580 2874.730 1074.590 ;
        RECT 2874.350 962.690 2874.730 962.700 ;
        RECT 2917.600 962.690 2924.800 963.140 ;
        RECT 2874.350 962.390 2924.800 962.690 ;
        RECT 2874.350 962.380 2874.730 962.390 ;
        RECT 2917.600 961.940 2924.800 962.390 ;
      LAYER met4 ;
        RECT 2874.375 1074.575 2874.705 1074.905 ;
        RECT 2874.390 962.705 2874.690 1074.575 ;
        RECT 2874.375 962.375 2874.705 962.705 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 1291.130 2873.810 1291.140 ;
        RECT 2859.820 1290.830 2873.810 1291.130 ;
        RECT 2873.430 1290.820 2873.810 1290.830 ;
        RECT 2873.430 1161.930 2873.810 1161.940 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2873.430 1161.630 2924.800 1161.930 ;
        RECT 2873.430 1161.620 2873.810 1161.630 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
      LAYER met4 ;
        RECT 2873.455 1290.815 2873.785 1291.145 ;
        RECT 2873.470 1161.945 2873.770 1290.815 ;
        RECT 2873.455 1161.615 2873.785 1161.945 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 1507.370 2873.810 1507.380 ;
        RECT 2859.820 1507.070 2873.810 1507.370 ;
        RECT 2873.430 1507.060 2873.810 1507.070 ;
        RECT 2873.430 1361.170 2873.810 1361.180 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2873.430 1360.870 2924.800 1361.170 ;
        RECT 2873.430 1360.860 2873.810 1360.870 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
      LAYER met4 ;
        RECT 2873.455 1507.055 2873.785 1507.385 ;
        RECT 2873.470 1361.185 2873.770 1507.055 ;
        RECT 2873.455 1360.855 2873.785 1361.185 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 1723.610 2873.810 1723.620 ;
        RECT 2859.820 1723.310 2873.810 1723.610 ;
        RECT 2873.430 1723.300 2873.810 1723.310 ;
        RECT 2873.430 1626.370 2873.810 1626.380 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2873.430 1626.070 2924.800 1626.370 ;
        RECT 2873.430 1626.060 2873.810 1626.070 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
      LAYER met4 ;
        RECT 2873.455 1723.295 2873.785 1723.625 ;
        RECT 2873.470 1626.385 2873.770 1723.295 ;
        RECT 2873.455 1626.055 2873.785 1626.385 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2877.110 137.850 2877.490 137.860 ;
        RECT 2859.820 137.550 2877.490 137.850 ;
        RECT 2877.110 137.540 2877.490 137.550 ;
        RECT 2877.110 99.090 2877.490 99.100 ;
        RECT 2917.600 99.090 2924.800 99.540 ;
        RECT 2877.110 98.790 2924.800 99.090 ;
        RECT 2877.110 98.780 2877.490 98.790 ;
        RECT 2917.600 98.340 2924.800 98.790 ;
      LAYER met4 ;
        RECT 2877.135 137.535 2877.465 137.865 ;
        RECT 2877.150 99.105 2877.450 137.535 ;
        RECT 2877.135 98.775 2877.465 99.105 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 354.090 2873.810 354.100 ;
        RECT 2859.820 353.790 2873.810 354.090 ;
        RECT 2873.430 353.780 2873.810 353.790 ;
        RECT 2873.430 298.330 2873.810 298.340 ;
        RECT 2917.600 298.330 2924.800 298.780 ;
        RECT 2873.430 298.030 2924.800 298.330 ;
        RECT 2873.430 298.020 2873.810 298.030 ;
        RECT 2917.600 297.580 2924.800 298.030 ;
      LAYER met4 ;
        RECT 2873.455 353.775 2873.785 354.105 ;
        RECT 2873.470 298.345 2873.770 353.775 ;
        RECT 2873.455 298.015 2873.785 298.345 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 570.330 2873.810 570.340 ;
        RECT 2859.820 570.030 2873.810 570.330 ;
        RECT 2873.430 570.020 2873.810 570.030 ;
        RECT 2873.430 497.570 2873.810 497.580 ;
        RECT 2917.600 497.570 2924.800 498.020 ;
        RECT 2873.430 497.270 2924.800 497.570 ;
        RECT 2873.430 497.260 2873.810 497.270 ;
        RECT 2917.600 496.820 2924.800 497.270 ;
      LAYER met4 ;
        RECT 2873.455 570.015 2873.785 570.345 ;
        RECT 2873.470 497.585 2873.770 570.015 ;
        RECT 2873.455 497.255 2873.785 497.585 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1792.290 2.400 1792.740 ;
        RECT 17.750 1792.290 18.130 1792.300 ;
        RECT -4.800 1791.990 18.130 1792.290 ;
        RECT -4.800 1791.540 2.400 1791.990 ;
        RECT 17.750 1791.980 18.130 1791.990 ;
        RECT 17.750 1651.530 18.130 1651.540 ;
        RECT 17.750 1651.230 60.260 1651.530 ;
        RECT 17.750 1651.220 18.130 1651.230 ;
      LAYER met4 ;
        RECT 17.775 1791.975 18.105 1792.305 ;
        RECT 17.790 1651.545 18.090 1791.975 ;
        RECT 17.775 1651.215 18.105 1651.545 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1531.170 2.400 1531.620 ;
        RECT 17.750 1531.170 18.130 1531.180 ;
        RECT -4.800 1530.870 18.130 1531.170 ;
        RECT -4.800 1530.420 2.400 1530.870 ;
        RECT 17.750 1530.860 18.130 1530.870 ;
        RECT 17.750 1435.290 18.130 1435.300 ;
        RECT 17.750 1434.990 60.260 1435.290 ;
        RECT 17.750 1434.980 18.130 1434.990 ;
      LAYER met4 ;
        RECT 17.775 1530.855 18.105 1531.185 ;
        RECT 17.790 1435.305 18.090 1530.855 ;
        RECT 17.775 1434.975 18.105 1435.305 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1270.730 2.400 1271.180 ;
        RECT 37.070 1270.730 37.450 1270.740 ;
        RECT -4.800 1270.430 37.450 1270.730 ;
        RECT -4.800 1269.980 2.400 1270.430 ;
        RECT 37.070 1270.420 37.450 1270.430 ;
        RECT 37.070 1219.050 37.450 1219.060 ;
        RECT 37.070 1218.750 60.260 1219.050 ;
        RECT 37.070 1218.740 37.450 1218.750 ;
      LAYER met4 ;
        RECT 37.095 1270.415 37.425 1270.745 ;
        RECT 37.110 1219.065 37.410 1270.415 ;
        RECT 37.095 1218.735 37.425 1219.065 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1009.610 2.400 1010.060 ;
        RECT -4.800 1009.310 34.650 1009.610 ;
        RECT -4.800 1008.860 2.400 1009.310 ;
        RECT 34.350 1006.210 34.650 1009.310 ;
        RECT 34.350 1005.910 60.410 1006.210 ;
        RECT 60.110 1002.660 60.410 1005.910 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.550 786.570 31.930 786.580 ;
        RECT 31.550 786.270 60.260 786.570 ;
        RECT 31.550 786.260 31.930 786.270 ;
        RECT -4.800 749.170 2.400 749.620 ;
        RECT 31.550 749.170 31.930 749.180 ;
        RECT -4.800 748.870 31.930 749.170 ;
        RECT -4.800 748.420 2.400 748.870 ;
        RECT 31.550 748.860 31.930 748.870 ;
      LAYER met4 ;
        RECT 31.575 786.255 31.905 786.585 ;
        RECT 31.590 749.185 31.890 786.255 ;
        RECT 31.575 748.855 31.905 749.185 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.750 570.330 18.130 570.340 ;
        RECT 17.750 570.030 60.260 570.330 ;
        RECT 17.750 570.020 18.130 570.030 ;
        RECT -4.800 488.050 2.400 488.500 ;
        RECT 17.750 488.050 18.130 488.060 ;
        RECT -4.800 487.750 18.130 488.050 ;
        RECT -4.800 487.300 2.400 487.750 ;
        RECT 17.750 487.740 18.130 487.750 ;
      LAYER met4 ;
        RECT 17.775 570.015 18.105 570.345 ;
        RECT 17.790 488.065 18.090 570.015 ;
        RECT 17.775 487.735 18.105 488.065 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.430 354.090 44.810 354.100 ;
        RECT 44.430 353.790 60.260 354.090 ;
        RECT 44.430 353.780 44.810 353.790 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 44.430 292.890 44.810 292.900 ;
        RECT -4.800 292.590 44.810 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 44.430 292.580 44.810 292.590 ;
      LAYER met4 ;
        RECT 44.455 353.775 44.785 354.105 ;
        RECT 44.470 292.905 44.770 353.775 ;
        RECT 44.455 292.575 44.785 292.905 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.550 137.850 31.930 137.860 ;
        RECT 31.550 137.550 60.260 137.850 ;
        RECT 31.550 137.540 31.930 137.550 ;
        RECT -4.800 97.050 2.400 97.500 ;
        RECT 31.550 97.050 31.930 97.060 ;
        RECT -4.800 96.750 31.930 97.050 ;
        RECT -4.800 96.300 2.400 96.750 ;
        RECT 31.550 96.740 31.930 96.750 ;
      LAYER met4 ;
        RECT 31.575 137.535 31.905 137.865 ;
        RECT 31.590 97.065 31.890 137.535 ;
        RECT 31.575 96.735 31.905 97.065 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 786.570 2874.730 786.580 ;
        RECT 2859.820 786.270 2874.730 786.570 ;
        RECT 2874.350 786.260 2874.730 786.270 ;
        RECT 2874.350 696.810 2874.730 696.820 ;
        RECT 2917.600 696.810 2924.800 697.260 ;
        RECT 2874.350 696.510 2924.800 696.810 ;
        RECT 2874.350 696.500 2874.730 696.510 ;
        RECT 2917.600 696.060 2924.800 696.510 ;
      LAYER met4 ;
        RECT 2874.375 786.255 2874.705 786.585 ;
        RECT 2874.390 696.825 2874.690 786.255 ;
        RECT 2874.375 696.495 2874.705 696.825 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2873.430 1002.810 2873.810 1002.820 ;
        RECT 2859.820 1002.510 2873.810 1002.810 ;
        RECT 2873.430 1002.500 2873.810 1002.510 ;
        RECT 2873.430 896.050 2873.810 896.060 ;
        RECT 2917.600 896.050 2924.800 896.500 ;
        RECT 2873.430 895.750 2924.800 896.050 ;
        RECT 2873.430 895.740 2873.810 895.750 ;
        RECT 2917.600 895.300 2924.800 895.750 ;
      LAYER met4 ;
        RECT 2873.455 1002.495 2873.785 1002.825 ;
        RECT 2873.470 896.065 2873.770 1002.495 ;
        RECT 2873.455 895.735 2873.785 896.065 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 1219.050 2874.730 1219.060 ;
        RECT 2859.820 1218.750 2874.730 1219.050 ;
        RECT 2874.350 1218.740 2874.730 1218.750 ;
        RECT 2874.350 1095.290 2874.730 1095.300 ;
        RECT 2917.600 1095.290 2924.800 1095.740 ;
        RECT 2874.350 1094.990 2924.800 1095.290 ;
        RECT 2874.350 1094.980 2874.730 1094.990 ;
        RECT 2917.600 1094.540 2924.800 1094.990 ;
      LAYER met4 ;
        RECT 2874.375 1218.735 2874.705 1219.065 ;
        RECT 2874.390 1095.305 2874.690 1218.735 ;
        RECT 2874.375 1094.975 2874.705 1095.305 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2875.270 1435.290 2875.650 1435.300 ;
        RECT 2859.820 1434.990 2875.650 1435.290 ;
        RECT 2875.270 1434.980 2875.650 1434.990 ;
        RECT 2875.270 1294.530 2875.650 1294.540 ;
        RECT 2917.600 1294.530 2924.800 1294.980 ;
        RECT 2875.270 1294.230 2924.800 1294.530 ;
        RECT 2875.270 1294.220 2875.650 1294.230 ;
        RECT 2917.600 1293.780 2924.800 1294.230 ;
      LAYER met4 ;
        RECT 2875.295 1434.975 2875.625 1435.305 ;
        RECT 2875.310 1294.545 2875.610 1434.975 ;
        RECT 2875.295 1294.215 2875.625 1294.545 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2874.350 1651.530 2874.730 1651.540 ;
        RECT 2859.820 1651.230 2874.730 1651.530 ;
        RECT 2874.350 1651.220 2874.730 1651.230 ;
        RECT 2874.350 1560.410 2874.730 1560.420 ;
        RECT 2917.600 1560.410 2924.800 1560.860 ;
        RECT 2874.350 1560.110 2924.800 1560.410 ;
        RECT 2874.350 1560.100 2874.730 1560.110 ;
        RECT 2917.600 1559.660 2924.800 1560.110 ;
      LAYER met4 ;
        RECT 2874.375 1651.215 2874.705 1651.545 ;
        RECT 2874.390 1560.425 2874.690 1651.215 ;
        RECT 2874.375 1560.095 2874.705 1560.425 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.170 14.010 687.310 15.300 ;
        RECT 686.480 13.870 687.310 14.010 ;
        RECT 628.450 1.090 628.730 1.205 ;
        RECT 629.230 1.090 629.790 2.400 ;
        RECT 686.480 1.205 686.620 13.870 ;
        RECT 628.450 0.950 629.790 1.090 ;
        RECT 628.450 0.835 628.730 0.950 ;
        RECT 629.230 -4.800 629.790 0.950 ;
        RECT 686.410 0.835 686.690 1.205 ;
      LAYER met3 ;
        RECT 628.425 1.170 628.755 1.185 ;
        RECT 686.385 1.170 686.715 1.185 ;
        RECT 628.425 0.870 686.715 1.170 ;
        RECT 628.425 0.855 628.755 0.870 ;
        RECT 686.385 0.855 686.715 0.870 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.170 14.010 2343.310 15.300 ;
        RECT 2343.170 13.870 2343.540 14.010 ;
        RECT 2343.400 10.725 2343.540 13.870 ;
        RECT 2343.330 10.355 2343.610 10.725 ;
        RECT 2402.670 10.355 2402.950 10.725 ;
        RECT 2402.740 2.400 2402.880 10.355 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
      LAYER met3 ;
        RECT 2343.305 10.690 2343.635 10.705 ;
        RECT 2402.645 10.690 2402.975 10.705 ;
        RECT 2343.305 10.390 2402.975 10.690 ;
        RECT 2343.305 10.375 2343.635 10.390 ;
        RECT 2402.645 10.375 2402.975 10.390 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.730 14.805 2359.870 15.300 ;
        RECT 2359.660 14.435 2359.940 14.805 ;
        RECT 2419.690 13.755 2419.970 14.125 ;
        RECT 2419.760 9.930 2419.900 13.755 ;
        RECT 2419.760 9.790 2420.360 9.930 ;
        RECT 2420.220 2.400 2420.360 9.790 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
      LAYER met3 ;
        RECT 2359.635 14.770 2359.965 14.785 ;
        RECT 2359.635 14.470 2419.290 14.770 ;
        RECT 2359.635 14.455 2359.965 14.470 ;
        RECT 2418.990 14.090 2419.290 14.470 ;
        RECT 2419.665 14.090 2419.995 14.105 ;
        RECT 2418.990 13.790 2419.995 14.090 ;
        RECT 2419.665 13.775 2419.995 13.790 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.290 14.010 2376.430 15.300 ;
        RECT 2376.290 13.870 2376.660 14.010 ;
        RECT 2376.520 3.925 2376.660 13.870 ;
        RECT 2376.450 3.555 2376.730 3.925 ;
        RECT 2438.090 3.555 2438.370 3.925 ;
        RECT 2438.160 2.400 2438.300 3.555 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
      LAYER met3 ;
        RECT 2376.425 3.890 2376.755 3.905 ;
        RECT 2438.065 3.890 2438.395 3.905 ;
        RECT 2376.425 3.590 2438.395 3.890 ;
        RECT 2376.425 3.575 2376.755 3.590 ;
        RECT 2438.065 3.575 2438.395 3.590 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.850 14.010 2392.990 15.300 ;
        RECT 2392.850 13.870 2393.220 14.010 ;
        RECT 2393.080 2.565 2393.220 13.870 ;
        RECT 2393.010 2.195 2393.290 2.565 ;
        RECT 2453.730 2.195 2454.010 2.565 ;
        RECT 2453.800 1.770 2453.940 2.195 ;
        RECT 2455.430 1.770 2455.990 2.400 ;
        RECT 2453.800 1.630 2455.990 1.770 ;
        RECT 2455.430 -4.800 2455.990 1.630 ;
      LAYER met3 ;
        RECT 2392.985 2.530 2393.315 2.545 ;
        RECT 2453.705 2.530 2454.035 2.545 ;
        RECT 2392.985 2.230 2454.035 2.530 ;
        RECT 2392.985 2.215 2393.315 2.230 ;
        RECT 2453.705 2.215 2454.035 2.230 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2409.410 14.010 2409.550 15.300 ;
        RECT 2409.410 13.870 2409.780 14.010 ;
        RECT 2409.640 4.605 2409.780 13.870 ;
        RECT 2409.570 4.235 2409.850 4.605 ;
        RECT 2473.510 4.235 2473.790 4.605 ;
        RECT 2473.580 2.400 2473.720 4.235 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
      LAYER met3 ;
        RECT 2409.545 4.570 2409.875 4.585 ;
        RECT 2473.485 4.570 2473.815 4.585 ;
        RECT 2409.545 4.270 2473.815 4.570 ;
        RECT 2409.545 4.255 2409.875 4.270 ;
        RECT 2473.485 4.255 2473.815 4.270 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.970 14.805 2426.110 15.300 ;
        RECT 2425.900 14.435 2426.180 14.805 ;
        RECT 2490.990 12.395 2491.270 12.765 ;
        RECT 2491.060 2.400 2491.200 12.395 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
      LAYER met3 ;
        RECT 2490.710 15.450 2491.090 15.460 ;
        RECT 2449.350 15.150 2491.090 15.450 ;
        RECT 2425.875 14.770 2426.205 14.785 ;
        RECT 2449.350 14.770 2449.650 15.150 ;
        RECT 2490.710 15.140 2491.090 15.150 ;
        RECT 2425.875 14.470 2449.650 14.770 ;
        RECT 2425.875 14.455 2426.205 14.470 ;
        RECT 2490.965 12.740 2491.295 12.745 ;
        RECT 2490.710 12.730 2491.295 12.740 ;
        RECT 2490.710 12.430 2491.520 12.730 ;
        RECT 2490.710 12.420 2491.295 12.430 ;
        RECT 2490.965 12.415 2491.295 12.420 ;
      LAYER met4 ;
        RECT 2490.735 15.135 2491.065 15.465 ;
        RECT 2490.750 12.745 2491.050 15.135 ;
        RECT 2490.735 12.415 2491.065 12.745 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2442.210 6.360 2442.530 6.420 ;
        RECT 2508.450 6.360 2508.770 6.420 ;
        RECT 2442.210 6.220 2508.770 6.360 ;
        RECT 2442.210 6.160 2442.530 6.220 ;
        RECT 2508.450 6.160 2508.770 6.220 ;
      LAYER met2 ;
        RECT 2442.530 14.010 2442.670 15.300 ;
        RECT 2442.300 13.870 2442.670 14.010 ;
        RECT 2442.300 6.450 2442.440 13.870 ;
        RECT 2442.240 6.130 2442.500 6.450 ;
        RECT 2508.480 6.130 2508.740 6.450 ;
        RECT 2508.540 3.300 2508.680 6.130 ;
        RECT 2508.540 3.160 2509.140 3.300 ;
        RECT 2509.000 2.400 2509.140 3.160 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2459.090 14.125 2459.230 15.300 ;
        RECT 2459.020 13.755 2459.300 14.125 ;
        RECT 2526.870 13.755 2527.150 14.125 ;
        RECT 2526.940 2.400 2527.080 13.755 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
      LAYER met3 ;
        RECT 2458.995 14.090 2459.325 14.105 ;
        RECT 2526.845 14.090 2527.175 14.105 ;
        RECT 2458.995 13.790 2527.175 14.090 ;
        RECT 2458.995 13.775 2459.325 13.790 ;
        RECT 2526.845 13.775 2527.175 13.790 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2475.650 14.805 2475.790 15.300 ;
        RECT 2475.580 14.435 2475.860 14.805 ;
        RECT 2544.350 13.755 2544.630 14.125 ;
        RECT 2544.420 2.400 2544.560 13.755 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
      LAYER met3 ;
        RECT 2475.555 14.770 2475.885 14.785 ;
        RECT 2475.555 14.470 2540.730 14.770 ;
        RECT 2475.555 14.455 2475.885 14.470 ;
        RECT 2540.430 14.090 2540.730 14.470 ;
        RECT 2544.325 14.090 2544.655 14.105 ;
        RECT 2540.430 13.790 2544.655 14.090 ;
        RECT 2544.325 13.775 2544.655 13.790 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.210 14.010 2492.350 15.300 ;
        RECT 2492.210 13.870 2492.580 14.010 ;
        RECT 2492.440 3.245 2492.580 13.870 ;
        RECT 2492.370 2.875 2492.650 3.245 ;
        RECT 2562.290 2.875 2562.570 3.245 ;
        RECT 2562.360 2.400 2562.500 2.875 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
      LAYER met3 ;
        RECT 2492.345 3.210 2492.675 3.225 ;
        RECT 2562.265 3.210 2562.595 3.225 ;
        RECT 2492.345 2.910 2562.595 3.210 ;
        RECT 2492.345 2.895 2492.675 2.910 ;
        RECT 2562.265 2.895 2562.595 2.910 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.770 14.010 852.910 15.300 ;
        RECT 852.540 13.870 852.910 14.010 ;
        RECT 852.540 10.045 852.680 13.870 ;
        RECT 806.470 9.675 806.750 10.045 ;
        RECT 852.470 9.675 852.750 10.045 ;
        RECT 806.540 2.400 806.680 9.675 ;
        RECT 806.330 -4.800 806.890 2.400 ;
      LAYER met3 ;
        RECT 806.445 10.010 806.775 10.025 ;
        RECT 852.445 10.010 852.775 10.025 ;
        RECT 806.445 9.710 852.775 10.010 ;
        RECT 806.445 9.695 806.775 9.710 ;
        RECT 852.445 9.695 852.775 9.710 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.770 14.010 2508.910 15.300 ;
        RECT 2508.770 13.870 2510.520 14.010 ;
        RECT 2510.380 1.885 2510.520 13.870 ;
        RECT 2510.310 1.515 2510.590 1.885 ;
        RECT 2577.470 1.770 2577.750 1.885 ;
        RECT 2579.630 1.770 2580.190 2.400 ;
        RECT 2577.470 1.630 2580.190 1.770 ;
        RECT 2577.470 1.515 2577.750 1.630 ;
        RECT 2579.630 -4.800 2580.190 1.630 ;
      LAYER met3 ;
        RECT 2510.285 1.850 2510.615 1.865 ;
        RECT 2577.445 1.850 2577.775 1.865 ;
        RECT 2510.285 1.550 2577.775 1.850 ;
        RECT 2510.285 1.535 2510.615 1.550 ;
        RECT 2577.445 1.535 2577.775 1.550 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2525.010 1.260 2525.330 1.320 ;
        RECT 2598.610 1.260 2598.930 1.320 ;
        RECT 2525.010 1.120 2598.930 1.260 ;
        RECT 2525.010 1.060 2525.330 1.120 ;
        RECT 2598.610 1.060 2598.930 1.120 ;
      LAYER met2 ;
        RECT 2525.330 14.010 2525.470 15.300 ;
        RECT 2525.100 13.870 2525.470 14.010 ;
        RECT 2525.100 1.350 2525.240 13.870 ;
        RECT 2525.040 1.030 2525.300 1.350 ;
        RECT 2597.570 1.090 2598.130 2.400 ;
        RECT 2598.640 1.090 2598.900 1.350 ;
        RECT 2597.570 1.030 2598.900 1.090 ;
        RECT 2597.570 0.950 2598.840 1.030 ;
        RECT 2597.570 -4.800 2598.130 0.950 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.890 14.805 2542.030 15.300 ;
        RECT 2541.820 14.435 2542.100 14.805 ;
        RECT 2615.190 12.395 2615.470 12.765 ;
        RECT 2615.260 2.400 2615.400 12.395 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
      LAYER met3 ;
        RECT 2589.150 18.170 2589.530 18.180 ;
        RECT 2545.950 17.870 2589.530 18.170 ;
        RECT 2541.795 14.770 2542.125 14.785 ;
        RECT 2545.950 14.770 2546.250 17.870 ;
        RECT 2589.150 17.860 2589.530 17.870 ;
        RECT 2589.150 15.450 2589.530 15.460 ;
        RECT 2614.910 15.450 2615.290 15.460 ;
        RECT 2589.150 15.150 2615.290 15.450 ;
        RECT 2589.150 15.140 2589.530 15.150 ;
        RECT 2614.910 15.140 2615.290 15.150 ;
        RECT 2541.795 14.470 2546.250 14.770 ;
        RECT 2541.795 14.455 2542.125 14.470 ;
        RECT 2615.165 12.740 2615.495 12.745 ;
        RECT 2614.910 12.730 2615.495 12.740 ;
        RECT 2614.910 12.430 2615.720 12.730 ;
        RECT 2614.910 12.420 2615.495 12.430 ;
        RECT 2615.165 12.415 2615.495 12.420 ;
      LAYER met4 ;
        RECT 2589.175 17.855 2589.505 18.185 ;
        RECT 2589.190 15.465 2589.490 17.855 ;
        RECT 2589.175 15.135 2589.505 15.465 ;
        RECT 2614.935 15.135 2615.265 15.465 ;
        RECT 2614.950 12.745 2615.250 15.135 ;
        RECT 2614.935 12.415 2615.265 12.745 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2558.450 14.805 2558.590 15.300 ;
        RECT 2558.380 14.435 2558.660 14.805 ;
        RECT 2632.670 13.330 2632.950 13.445 ;
        RECT 2632.670 13.190 2633.340 13.330 ;
        RECT 2632.670 13.075 2632.950 13.190 ;
        RECT 2633.200 2.400 2633.340 13.190 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
      LAYER met3 ;
        RECT 2587.350 15.830 2622.150 16.130 ;
        RECT 2558.355 14.770 2558.685 14.785 ;
        RECT 2587.350 14.770 2587.650 15.830 ;
        RECT 2621.850 15.450 2622.150 15.830 ;
        RECT 2632.390 15.450 2632.770 15.460 ;
        RECT 2621.850 15.150 2632.770 15.450 ;
        RECT 2632.390 15.140 2632.770 15.150 ;
        RECT 2558.355 14.470 2573.850 14.770 ;
        RECT 2558.355 14.455 2558.685 14.470 ;
        RECT 2573.550 14.090 2573.850 14.470 ;
        RECT 2585.510 14.470 2587.650 14.770 ;
        RECT 2585.510 14.090 2585.810 14.470 ;
        RECT 2573.550 13.790 2585.810 14.090 ;
        RECT 2632.645 13.420 2632.975 13.425 ;
        RECT 2632.390 13.410 2632.975 13.420 ;
        RECT 2632.390 13.110 2633.200 13.410 ;
        RECT 2632.390 13.100 2632.975 13.110 ;
        RECT 2632.645 13.095 2632.975 13.100 ;
      LAYER met4 ;
        RECT 2632.415 15.135 2632.745 15.465 ;
        RECT 2632.430 13.425 2632.730 15.135 ;
        RECT 2632.415 13.095 2632.745 13.425 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.010 14.805 2575.150 15.300 ;
        RECT 2574.940 14.435 2575.220 14.805 ;
        RECT 2650.150 13.330 2650.430 13.445 ;
        RECT 2650.150 13.190 2650.820 13.330 ;
        RECT 2650.150 13.075 2650.430 13.190 ;
        RECT 2650.680 2.400 2650.820 13.190 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
      LAYER met3 ;
        RECT 2583.630 17.490 2584.010 17.500 ;
        RECT 2583.630 17.190 2650.210 17.490 ;
        RECT 2583.630 17.180 2584.010 17.190 ;
        RECT 2649.910 16.140 2650.210 17.190 ;
        RECT 2649.870 15.820 2650.250 16.140 ;
        RECT 2574.915 14.770 2575.245 14.785 ;
        RECT 2583.630 14.770 2584.010 14.780 ;
        RECT 2574.915 14.470 2584.010 14.770 ;
        RECT 2574.915 14.455 2575.245 14.470 ;
        RECT 2583.630 14.460 2584.010 14.470 ;
        RECT 2650.125 13.420 2650.455 13.425 ;
        RECT 2649.870 13.410 2650.455 13.420 ;
        RECT 2649.870 13.110 2650.680 13.410 ;
        RECT 2649.870 13.100 2650.455 13.110 ;
        RECT 2650.125 13.095 2650.455 13.100 ;
      LAYER met4 ;
        RECT 2583.655 17.175 2583.985 17.505 ;
        RECT 2583.670 14.785 2583.970 17.175 ;
        RECT 2649.895 15.815 2650.225 16.145 ;
        RECT 2583.655 14.455 2583.985 14.785 ;
        RECT 2649.910 13.425 2650.210 15.815 ;
        RECT 2649.895 13.095 2650.225 13.425 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.570 14.805 2591.710 15.300 ;
        RECT 2591.500 14.435 2591.780 14.805 ;
        RECT 2666.710 13.330 2666.990 13.445 ;
        RECT 2666.710 13.190 2668.760 13.330 ;
        RECT 2666.710 13.075 2666.990 13.190 ;
        RECT 2668.620 2.400 2668.760 13.190 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
      LAYER met3 ;
        RECT 2591.475 14.770 2591.805 14.785 ;
        RECT 2591.475 14.470 2622.150 14.770 ;
        RECT 2591.475 14.455 2591.805 14.470 ;
        RECT 2621.850 14.090 2622.150 14.470 ;
        RECT 2666.430 14.090 2666.810 14.100 ;
        RECT 2621.850 13.790 2666.810 14.090 ;
        RECT 2666.430 13.780 2666.810 13.790 ;
        RECT 2666.685 13.420 2667.015 13.425 ;
        RECT 2666.430 13.410 2667.015 13.420 ;
        RECT 2666.430 13.110 2667.240 13.410 ;
        RECT 2666.430 13.100 2667.015 13.110 ;
        RECT 2666.685 13.095 2667.015 13.100 ;
      LAYER met4 ;
        RECT 2666.455 13.775 2666.785 14.105 ;
        RECT 2666.470 13.425 2666.770 13.775 ;
        RECT 2666.455 13.095 2666.785 13.425 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2607.810 5.680 2608.130 5.740 ;
        RECT 2685.090 5.680 2685.410 5.740 ;
        RECT 2607.810 5.540 2685.410 5.680 ;
        RECT 2607.810 5.480 2608.130 5.540 ;
        RECT 2685.090 5.480 2685.410 5.540 ;
      LAYER met2 ;
        RECT 2608.130 14.010 2608.270 15.300 ;
        RECT 2607.900 13.870 2608.270 14.010 ;
        RECT 2607.900 5.770 2608.040 13.870 ;
        RECT 2685.180 5.770 2686.240 5.850 ;
        RECT 2607.840 5.450 2608.100 5.770 ;
        RECT 2685.120 5.710 2686.240 5.770 ;
        RECT 2685.120 5.450 2685.380 5.710 ;
        RECT 2686.100 2.400 2686.240 5.710 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2624.690 14.805 2624.830 15.300 ;
        RECT 2624.620 14.435 2624.900 14.805 ;
        RECT 2703.970 13.755 2704.250 14.125 ;
        RECT 2704.040 2.400 2704.180 13.755 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
      LAYER met3 ;
        RECT 2667.350 18.850 2667.730 18.860 ;
        RECT 2631.510 18.550 2667.730 18.850 ;
        RECT 2631.510 18.180 2631.810 18.550 ;
        RECT 2667.350 18.540 2667.730 18.550 ;
        RECT 2631.470 17.860 2631.850 18.180 ;
        RECT 2624.595 14.770 2624.925 14.785 ;
        RECT 2631.470 14.770 2631.850 14.780 ;
        RECT 2624.595 14.470 2631.850 14.770 ;
        RECT 2624.595 14.455 2624.925 14.470 ;
        RECT 2631.470 14.460 2631.850 14.470 ;
        RECT 2667.350 14.460 2667.730 14.780 ;
        RECT 2667.390 14.090 2667.690 14.460 ;
        RECT 2703.945 14.090 2704.275 14.105 ;
        RECT 2667.390 13.790 2704.275 14.090 ;
        RECT 2703.945 13.775 2704.275 13.790 ;
      LAYER met4 ;
        RECT 2667.375 18.535 2667.705 18.865 ;
        RECT 2631.495 17.855 2631.825 18.185 ;
        RECT 2631.510 14.785 2631.810 17.855 ;
        RECT 2667.390 14.785 2667.690 18.535 ;
        RECT 2631.495 14.455 2631.825 14.785 ;
        RECT 2667.375 14.455 2667.705 14.785 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2641.250 13.870 2641.390 15.300 ;
        RECT 2641.250 13.730 2641.620 13.870 ;
        RECT 2641.480 10.045 2641.620 13.730 ;
        RECT 2641.410 9.675 2641.690 10.045 ;
        RECT 2721.910 9.675 2722.190 10.045 ;
        RECT 2721.980 2.400 2722.120 9.675 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
      LAYER met3 ;
        RECT 2641.385 10.010 2641.715 10.025 ;
        RECT 2721.885 10.010 2722.215 10.025 ;
        RECT 2641.385 9.710 2722.215 10.010 ;
        RECT 2641.385 9.695 2641.715 9.710 ;
        RECT 2721.885 9.695 2722.215 9.710 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2657.810 14.805 2657.950 15.300 ;
        RECT 2657.740 14.435 2658.020 14.805 ;
        RECT 2739.390 12.395 2739.670 12.765 ;
        RECT 2739.460 2.400 2739.600 12.395 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
      LAYER met3 ;
        RECT 2738.190 17.490 2738.570 17.500 ;
        RECT 2674.750 17.190 2718.750 17.490 ;
        RECT 2666.700 15.150 2670.450 15.450 ;
        RECT 2657.715 14.770 2658.045 14.785 ;
        RECT 2666.700 14.770 2667.000 15.150 ;
        RECT 2657.715 14.470 2667.000 14.770 ;
        RECT 2670.150 14.770 2670.450 15.150 ;
        RECT 2674.750 14.770 2675.050 17.190 ;
        RECT 2718.450 16.810 2718.750 17.190 ;
        RECT 2727.190 17.190 2738.570 17.490 ;
        RECT 2727.190 16.810 2727.490 17.190 ;
        RECT 2738.190 17.180 2738.570 17.190 ;
        RECT 2718.450 16.510 2727.490 16.810 ;
        RECT 2670.150 14.470 2675.050 14.770 ;
        RECT 2657.715 14.455 2658.045 14.470 ;
        RECT 2738.190 12.730 2738.570 12.740 ;
        RECT 2739.365 12.730 2739.695 12.745 ;
        RECT 2738.190 12.430 2739.695 12.730 ;
        RECT 2738.190 12.420 2738.570 12.430 ;
        RECT 2739.365 12.415 2739.695 12.430 ;
      LAYER met4 ;
        RECT 2738.215 17.175 2738.545 17.505 ;
        RECT 2738.230 12.745 2738.530 17.175 ;
        RECT 2738.215 12.415 2738.545 12.745 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.330 14.010 869.470 15.300 ;
        RECT 869.100 13.870 869.470 14.010 ;
        RECT 869.100 6.645 869.240 13.870 ;
        RECT 824.410 6.275 824.690 6.645 ;
        RECT 869.030 6.275 869.310 6.645 ;
        RECT 824.480 2.400 824.620 6.275 ;
        RECT 824.270 -4.800 824.830 2.400 ;
      LAYER met3 ;
        RECT 824.385 6.610 824.715 6.625 ;
        RECT 869.005 6.610 869.335 6.625 ;
        RECT 824.385 6.310 869.335 6.610 ;
        RECT 824.385 6.295 824.715 6.310 ;
        RECT 869.005 6.295 869.335 6.310 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.370 14.010 2674.510 15.300 ;
        RECT 2674.370 13.870 2674.740 14.010 ;
        RECT 2674.600 3.925 2674.740 13.870 ;
        RECT 2674.530 3.555 2674.810 3.925 ;
        RECT 2757.400 2.990 2758.460 3.130 ;
        RECT 2757.400 2.400 2757.540 2.990 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
        RECT 2758.320 1.885 2758.460 2.990 ;
        RECT 2758.250 1.515 2758.530 1.885 ;
      LAYER met3 ;
        RECT 2674.505 3.890 2674.835 3.905 ;
        RECT 2674.505 3.590 2691.150 3.890 ;
        RECT 2674.505 3.575 2674.835 3.590 ;
        RECT 2690.850 1.850 2691.150 3.590 ;
        RECT 2758.225 1.850 2758.555 1.865 ;
        RECT 2690.850 1.550 2758.555 1.850 ;
        RECT 2758.225 1.535 2758.555 1.550 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2690.610 1.260 2690.930 1.320 ;
        RECT 2773.870 1.260 2774.190 1.320 ;
        RECT 2690.610 1.120 2774.190 1.260 ;
        RECT 2690.610 1.060 2690.930 1.120 ;
        RECT 2773.870 1.060 2774.190 1.120 ;
      LAYER met2 ;
        RECT 2690.930 14.010 2691.070 15.300 ;
        RECT 2690.700 13.870 2691.070 14.010 ;
        RECT 2690.700 1.350 2690.840 13.870 ;
        RECT 2690.640 1.030 2690.900 1.350 ;
        RECT 2773.900 1.090 2774.160 1.350 ;
        RECT 2774.670 1.090 2775.230 2.400 ;
        RECT 2773.900 1.030 2775.230 1.090 ;
        RECT 2773.960 0.950 2775.230 1.030 ;
        RECT 2774.670 -4.800 2775.230 0.950 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2707.490 14.805 2707.630 15.300 ;
        RECT 2707.420 14.435 2707.700 14.805 ;
        RECT 2792.750 13.755 2793.030 14.125 ;
        RECT 2792.820 2.400 2792.960 13.755 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
      LAYER met3 ;
        RECT 2792.470 19.530 2792.850 19.540 ;
        RECT 2766.750 19.230 2792.850 19.530 ;
        RECT 2766.750 16.130 2767.050 19.230 ;
        RECT 2792.470 19.220 2792.850 19.230 ;
        RECT 2739.150 15.830 2767.050 16.130 ;
        RECT 2707.395 14.770 2707.725 14.785 ;
        RECT 2739.150 14.770 2739.450 15.830 ;
        RECT 2707.395 14.470 2739.450 14.770 ;
        RECT 2707.395 14.455 2707.725 14.470 ;
        RECT 2792.725 14.100 2793.055 14.105 ;
        RECT 2792.470 14.090 2793.055 14.100 ;
        RECT 2792.470 13.790 2793.280 14.090 ;
        RECT 2792.470 13.780 2793.055 13.790 ;
        RECT 2792.725 13.775 2793.055 13.780 ;
      LAYER met4 ;
        RECT 2792.495 19.215 2792.825 19.545 ;
        RECT 2792.510 14.105 2792.810 19.215 ;
        RECT 2792.495 13.775 2792.825 14.105 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2724.050 13.870 2724.190 15.300 ;
        RECT 2724.050 13.730 2724.420 13.870 ;
        RECT 2724.280 0.525 2724.420 13.730 ;
        RECT 2724.210 0.155 2724.490 0.525 ;
        RECT 2810.090 0.410 2810.650 2.400 ;
        RECT 2811.150 0.410 2811.430 0.525 ;
        RECT 2810.090 0.270 2811.430 0.410 ;
        RECT 2810.090 -4.800 2810.650 0.270 ;
        RECT 2811.150 0.155 2811.430 0.270 ;
      LAYER met3 ;
        RECT 2724.185 0.490 2724.515 0.505 ;
        RECT 2811.125 0.490 2811.455 0.505 ;
        RECT 2724.185 0.190 2811.455 0.490 ;
        RECT 2724.185 0.175 2724.515 0.190 ;
        RECT 2811.125 0.175 2811.455 0.190 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2740.610 14.805 2740.750 15.300 ;
        RECT 2740.540 14.435 2740.820 14.805 ;
        RECT 2828.170 13.755 2828.450 14.125 ;
        RECT 2828.240 2.400 2828.380 13.755 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
      LAYER met3 ;
        RECT 2787.450 15.150 2810.290 15.450 ;
        RECT 2740.515 14.770 2740.845 14.785 ;
        RECT 2787.450 14.770 2787.750 15.150 ;
        RECT 2740.515 14.470 2787.750 14.770 ;
        RECT 2740.515 14.455 2740.845 14.470 ;
        RECT 2809.990 14.090 2810.290 15.150 ;
        RECT 2828.145 14.090 2828.475 14.105 ;
        RECT 2809.990 13.790 2828.475 14.090 ;
        RECT 2828.145 13.775 2828.475 13.790 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.170 13.870 2757.310 15.300 ;
        RECT 2756.940 13.730 2757.310 13.870 ;
        RECT 2756.940 3.245 2757.080 13.730 ;
        RECT 2756.870 2.875 2757.150 3.245 ;
        RECT 2845.650 2.875 2845.930 3.245 ;
        RECT 2845.720 2.400 2845.860 2.875 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
      LAYER met3 ;
        RECT 2756.845 3.210 2757.175 3.225 ;
        RECT 2845.625 3.210 2845.955 3.225 ;
        RECT 2756.845 2.910 2845.955 3.210 ;
        RECT 2756.845 2.895 2757.175 2.910 ;
        RECT 2845.625 2.895 2845.955 2.910 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2773.410 1.600 2773.730 1.660 ;
        RECT 2864.490 1.600 2864.810 1.660 ;
        RECT 2773.410 1.460 2864.810 1.600 ;
        RECT 2773.410 1.400 2773.730 1.460 ;
        RECT 2864.490 1.400 2864.810 1.460 ;
      LAYER met2 ;
        RECT 2773.730 14.010 2773.870 15.300 ;
        RECT 2773.500 13.870 2773.870 14.010 ;
        RECT 2773.500 1.690 2773.640 13.870 ;
        RECT 2863.450 1.770 2864.010 2.400 ;
        RECT 2863.450 1.690 2864.720 1.770 ;
        RECT 2773.440 1.370 2773.700 1.690 ;
        RECT 2863.450 1.630 2864.780 1.690 ;
        RECT 2863.450 -4.800 2864.010 1.630 ;
        RECT 2864.520 1.370 2864.780 1.630 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2790.290 14.010 2790.430 15.300 ;
        RECT 2790.290 13.870 2790.660 14.010 ;
        RECT 2790.520 1.885 2790.660 13.870 ;
        RECT 2790.450 1.515 2790.730 1.885 ;
        RECT 2878.770 1.770 2879.050 1.885 ;
        RECT 2881.390 1.770 2881.950 2.400 ;
        RECT 2878.770 1.630 2881.950 1.770 ;
        RECT 2878.770 1.515 2879.050 1.630 ;
        RECT 2881.390 -4.800 2881.950 1.630 ;
      LAYER met3 ;
        RECT 2790.425 1.850 2790.755 1.865 ;
        RECT 2878.745 1.850 2879.075 1.865 ;
        RECT 2790.425 1.550 2879.075 1.850 ;
        RECT 2790.425 1.535 2790.755 1.550 ;
        RECT 2878.745 1.535 2879.075 1.550 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.890 14.010 886.030 15.300 ;
        RECT 885.660 13.870 886.030 14.010 ;
        RECT 885.660 5.285 885.800 13.870 ;
        RECT 841.890 4.915 842.170 5.285 ;
        RECT 885.590 4.915 885.870 5.285 ;
        RECT 841.960 2.400 842.100 4.915 ;
        RECT 841.750 -4.800 842.310 2.400 ;
      LAYER met3 ;
        RECT 841.865 5.250 842.195 5.265 ;
        RECT 885.565 5.250 885.895 5.265 ;
        RECT 841.865 4.950 885.895 5.250 ;
        RECT 841.865 4.935 842.195 4.950 ;
        RECT 885.565 4.935 885.895 4.950 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.450 14.010 902.590 15.300 ;
        RECT 902.220 13.870 902.590 14.010 ;
        RECT 902.220 5.965 902.360 13.870 ;
        RECT 859.830 5.595 860.110 5.965 ;
        RECT 902.150 5.595 902.430 5.965 ;
        RECT 859.900 2.400 860.040 5.595 ;
        RECT 859.690 -4.800 860.250 2.400 ;
      LAYER met3 ;
        RECT 859.805 5.930 860.135 5.945 ;
        RECT 902.125 5.930 902.455 5.945 ;
        RECT 859.805 5.630 902.455 5.930 ;
        RECT 859.805 5.615 860.135 5.630 ;
        RECT 902.125 5.615 902.455 5.630 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.010 14.010 919.150 15.300 ;
        RECT 917.860 13.870 919.150 14.010 ;
        RECT 877.170 0.410 877.730 2.400 ;
        RECT 879.150 0.410 879.430 0.525 ;
        RECT 877.170 0.270 879.430 0.410 ;
        RECT 877.170 -4.800 877.730 0.270 ;
        RECT 879.150 0.155 879.430 0.270 ;
        RECT 917.330 0.410 917.610 0.525 ;
        RECT 917.860 0.410 918.000 13.870 ;
        RECT 917.330 0.270 918.000 0.410 ;
        RECT 917.330 0.155 917.610 0.270 ;
      LAYER met3 ;
        RECT 879.125 0.490 879.455 0.505 ;
        RECT 917.305 0.490 917.635 0.505 ;
        RECT 879.125 0.190 917.635 0.490 ;
        RECT 879.125 0.175 879.455 0.190 ;
        RECT 917.305 0.175 917.635 0.190 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.570 14.010 935.710 15.300 ;
        RECT 935.340 13.870 935.710 14.010 ;
        RECT 935.340 3.925 935.480 13.870 ;
        RECT 895.250 3.555 895.530 3.925 ;
        RECT 935.270 3.555 935.550 3.925 ;
        RECT 895.320 2.400 895.460 3.555 ;
        RECT 895.110 -4.800 895.670 2.400 ;
      LAYER met3 ;
        RECT 895.225 3.890 895.555 3.905 ;
        RECT 935.245 3.890 935.575 3.905 ;
        RECT 895.225 3.590 935.575 3.890 ;
        RECT 895.225 3.575 895.555 3.590 ;
        RECT 935.245 3.575 935.575 3.590 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.130 14.010 952.270 15.300 ;
        RECT 951.900 13.870 952.270 14.010 ;
        RECT 911.810 1.090 912.090 1.205 ;
        RECT 912.590 1.090 913.150 2.400 ;
        RECT 951.900 1.205 952.040 13.870 ;
        RECT 911.810 0.950 913.150 1.090 ;
        RECT 911.810 0.835 912.090 0.950 ;
        RECT 912.590 -4.800 913.150 0.950 ;
        RECT 951.830 0.835 952.110 1.205 ;
      LAYER met3 ;
        RECT 911.785 1.170 912.115 1.185 ;
        RECT 951.805 1.170 952.135 1.185 ;
        RECT 911.785 0.870 952.135 1.170 ;
        RECT 911.785 0.855 912.115 0.870 ;
        RECT 951.805 0.855 952.135 0.870 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.690 14.125 968.830 15.300 ;
        RECT 930.670 13.755 930.950 14.125 ;
        RECT 968.620 13.755 968.900 14.125 ;
        RECT 930.740 2.400 930.880 13.755 ;
        RECT 930.530 -4.800 931.090 2.400 ;
      LAYER met3 ;
        RECT 930.645 14.090 930.975 14.105 ;
        RECT 968.595 14.090 968.925 14.105 ;
        RECT 930.645 13.790 968.925 14.090 ;
        RECT 930.645 13.775 930.975 13.790 ;
        RECT 968.595 13.775 968.925 13.790 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.250 14.010 985.390 15.300 ;
        RECT 985.020 13.870 985.390 14.010 ;
        RECT 985.020 10.045 985.160 13.870 ;
        RECT 948.610 9.675 948.890 10.045 ;
        RECT 984.950 9.675 985.230 10.045 ;
        RECT 948.680 2.400 948.820 9.675 ;
        RECT 948.470 -4.800 949.030 2.400 ;
      LAYER met3 ;
        RECT 948.585 10.010 948.915 10.025 ;
        RECT 984.925 10.010 985.255 10.025 ;
        RECT 948.585 9.710 985.255 10.010 ;
        RECT 948.585 9.695 948.915 9.710 ;
        RECT 984.925 9.695 985.255 9.710 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.810 14.010 1001.950 15.300 ;
        RECT 1001.580 13.870 1001.950 14.010 ;
        RECT 1001.580 5.285 1001.720 13.870 ;
        RECT 966.090 4.915 966.370 5.285 ;
        RECT 1001.510 4.915 1001.790 5.285 ;
        RECT 966.160 2.400 966.300 4.915 ;
        RECT 965.950 -4.800 966.510 2.400 ;
      LAYER met3 ;
        RECT 966.065 5.250 966.395 5.265 ;
        RECT 1001.485 5.250 1001.815 5.265 ;
        RECT 966.065 4.950 1001.815 5.250 ;
        RECT 966.065 4.935 966.395 4.950 ;
        RECT 1001.485 4.935 1001.815 4.950 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.730 14.010 703.870 15.300 ;
        RECT 703.500 13.870 703.870 14.010 ;
        RECT 703.500 4.605 703.640 13.870 ;
        RECT 646.850 4.235 647.130 4.605 ;
        RECT 703.430 4.235 703.710 4.605 ;
        RECT 646.920 2.400 647.060 4.235 ;
        RECT 646.710 -4.800 647.270 2.400 ;
      LAYER met3 ;
        RECT 646.825 4.570 647.155 4.585 ;
        RECT 703.405 4.570 703.735 4.585 ;
        RECT 646.825 4.270 703.735 4.570 ;
        RECT 646.825 4.255 647.155 4.270 ;
        RECT 703.405 4.255 703.735 4.270 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.370 14.010 1018.510 15.300 ;
        RECT 1017.680 13.870 1018.510 14.010 ;
        RECT 983.890 0.410 984.450 2.400 ;
        RECT 1017.680 0.525 1017.820 13.870 ;
        RECT 985.870 0.410 986.150 0.525 ;
        RECT 983.890 0.270 986.150 0.410 ;
        RECT 983.890 -4.800 984.450 0.270 ;
        RECT 985.870 0.155 986.150 0.270 ;
        RECT 1017.610 0.155 1017.890 0.525 ;
      LAYER met3 ;
        RECT 985.845 0.490 986.175 0.505 ;
        RECT 1017.585 0.490 1017.915 0.505 ;
        RECT 985.845 0.190 1017.915 0.490 ;
        RECT 985.845 0.175 986.175 0.190 ;
        RECT 1017.585 0.175 1017.915 0.190 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.930 14.010 1035.070 15.300 ;
        RECT 1034.700 13.870 1035.070 14.010 ;
        RECT 1034.700 8.685 1034.840 13.870 ;
        RECT 1002.430 8.570 1002.710 8.685 ;
        RECT 1002.040 8.430 1002.710 8.570 ;
        RECT 1002.040 4.490 1002.180 8.430 ;
        RECT 1002.430 8.315 1002.710 8.430 ;
        RECT 1034.630 8.315 1034.910 8.685 ;
        RECT 1001.580 4.350 1002.180 4.490 ;
        RECT 1001.580 2.400 1001.720 4.350 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
      LAYER met3 ;
        RECT 1002.405 8.650 1002.735 8.665 ;
        RECT 1034.605 8.650 1034.935 8.665 ;
        RECT 1002.405 8.350 1034.935 8.650 ;
        RECT 1002.405 8.335 1002.735 8.350 ;
        RECT 1034.605 8.335 1034.935 8.350 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.490 14.010 1051.630 15.300 ;
        RECT 1051.260 13.870 1051.630 14.010 ;
        RECT 1051.260 5.965 1051.400 13.870 ;
        RECT 1019.450 5.595 1019.730 5.965 ;
        RECT 1051.190 5.595 1051.470 5.965 ;
        RECT 1019.520 2.400 1019.660 5.595 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER met3 ;
        RECT 1019.425 5.930 1019.755 5.945 ;
        RECT 1051.165 5.930 1051.495 5.945 ;
        RECT 1019.425 5.630 1051.495 5.930 ;
        RECT 1019.425 5.615 1019.755 5.630 ;
        RECT 1051.165 5.615 1051.495 5.630 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.050 14.010 1068.190 15.300 ;
        RECT 1067.820 13.870 1068.190 14.010 ;
        RECT 1067.820 10.725 1067.960 13.870 ;
        RECT 1036.930 10.355 1037.210 10.725 ;
        RECT 1067.750 10.355 1068.030 10.725 ;
        RECT 1037.000 2.400 1037.140 10.355 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
      LAYER met3 ;
        RECT 1036.905 10.690 1037.235 10.705 ;
        RECT 1067.725 10.690 1068.055 10.705 ;
        RECT 1036.905 10.390 1068.055 10.690 ;
        RECT 1036.905 10.375 1037.235 10.390 ;
        RECT 1067.725 10.375 1068.055 10.390 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.610 14.010 1084.750 15.300 ;
        RECT 1084.610 13.870 1084.980 14.010 ;
        RECT 1084.840 5.965 1084.980 13.870 ;
        RECT 1054.870 5.595 1055.150 5.965 ;
        RECT 1084.770 5.595 1085.050 5.965 ;
        RECT 1054.940 2.400 1055.080 5.595 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
      LAYER met3 ;
        RECT 1054.845 5.930 1055.175 5.945 ;
        RECT 1084.745 5.930 1085.075 5.945 ;
        RECT 1054.845 5.630 1085.075 5.930 ;
        RECT 1054.845 5.615 1055.175 5.630 ;
        RECT 1084.745 5.615 1085.075 5.630 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.170 14.010 1101.310 15.300 ;
        RECT 1100.940 13.870 1101.310 14.010 ;
        RECT 1100.940 7.325 1101.080 13.870 ;
        RECT 1072.350 6.955 1072.630 7.325 ;
        RECT 1100.870 6.955 1101.150 7.325 ;
        RECT 1072.420 2.400 1072.560 6.955 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
      LAYER met3 ;
        RECT 1072.325 7.290 1072.655 7.305 ;
        RECT 1100.845 7.290 1101.175 7.305 ;
        RECT 1072.325 6.990 1101.175 7.290 ;
        RECT 1072.325 6.975 1072.655 6.990 ;
        RECT 1100.845 6.975 1101.175 6.990 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.730 14.010 1117.870 15.300 ;
        RECT 1117.500 13.870 1117.870 14.010 ;
        RECT 1117.500 13.445 1117.640 13.870 ;
        RECT 1090.290 13.075 1090.570 13.445 ;
        RECT 1117.430 13.075 1117.710 13.445 ;
        RECT 1090.360 2.400 1090.500 13.075 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
      LAYER met3 ;
        RECT 1090.265 13.410 1090.595 13.425 ;
        RECT 1117.405 13.410 1117.735 13.425 ;
        RECT 1090.265 13.110 1117.735 13.410 ;
        RECT 1090.265 13.095 1090.595 13.110 ;
        RECT 1117.405 13.095 1117.735 13.110 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.290 14.010 1134.430 15.300 ;
        RECT 1134.060 13.870 1134.430 14.010 ;
        RECT 1134.060 9.365 1134.200 13.870 ;
        RECT 1107.770 8.995 1108.050 9.365 ;
        RECT 1133.990 8.995 1134.270 9.365 ;
        RECT 1107.840 2.400 1107.980 8.995 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
      LAYER met3 ;
        RECT 1107.745 9.330 1108.075 9.345 ;
        RECT 1133.965 9.330 1134.295 9.345 ;
        RECT 1107.745 9.030 1134.295 9.330 ;
        RECT 1107.745 9.015 1108.075 9.030 ;
        RECT 1133.965 9.015 1134.295 9.030 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.850 14.010 1150.990 15.300 ;
        RECT 1150.620 13.870 1150.990 14.010 ;
        RECT 1150.620 7.325 1150.760 13.870 ;
        RECT 1125.710 6.955 1125.990 7.325 ;
        RECT 1150.550 6.955 1150.830 7.325 ;
        RECT 1125.780 2.400 1125.920 6.955 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
      LAYER met3 ;
        RECT 1125.685 7.290 1126.015 7.305 ;
        RECT 1150.525 7.290 1150.855 7.305 ;
        RECT 1125.685 6.990 1150.855 7.290 ;
        RECT 1125.685 6.975 1126.015 6.990 ;
        RECT 1150.525 6.975 1150.855 6.990 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.410 14.010 1167.550 15.300 ;
        RECT 1167.180 13.870 1167.550 14.010 ;
        RECT 1167.180 12.085 1167.320 13.870 ;
        RECT 1143.650 11.715 1143.930 12.085 ;
        RECT 1167.110 11.715 1167.390 12.085 ;
        RECT 1143.720 2.400 1143.860 11.715 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
      LAYER met3 ;
        RECT 1143.625 12.050 1143.955 12.065 ;
        RECT 1167.085 12.050 1167.415 12.065 ;
        RECT 1143.625 11.750 1167.415 12.050 ;
        RECT 1143.625 11.735 1143.955 11.750 ;
        RECT 1167.085 11.735 1167.415 11.750 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.290 14.010 720.430 15.300 ;
        RECT 720.060 13.870 720.430 14.010 ;
        RECT 720.060 3.245 720.200 13.870 ;
        RECT 664.790 2.875 665.070 3.245 ;
        RECT 719.990 2.875 720.270 3.245 ;
        RECT 664.860 2.400 665.000 2.875 ;
        RECT 664.650 -4.800 665.210 2.400 ;
      LAYER met3 ;
        RECT 664.765 3.210 665.095 3.225 ;
        RECT 719.965 3.210 720.295 3.225 ;
        RECT 664.765 2.910 720.295 3.210 ;
        RECT 664.765 2.895 665.095 2.910 ;
        RECT 719.965 2.895 720.295 2.910 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.970 14.010 1184.110 15.300 ;
        RECT 1183.740 13.870 1184.110 14.010 ;
        RECT 1183.740 8.005 1183.880 13.870 ;
        RECT 1161.130 7.635 1161.410 8.005 ;
        RECT 1183.670 7.635 1183.950 8.005 ;
        RECT 1161.200 2.400 1161.340 7.635 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
      LAYER met3 ;
        RECT 1161.105 7.970 1161.435 7.985 ;
        RECT 1183.645 7.970 1183.975 7.985 ;
        RECT 1161.105 7.670 1183.975 7.970 ;
        RECT 1161.105 7.655 1161.435 7.670 ;
        RECT 1183.645 7.655 1183.975 7.670 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.530 14.010 1200.670 15.300 ;
        RECT 1200.300 13.870 1200.670 14.010 ;
        RECT 1200.300 7.325 1200.440 13.870 ;
        RECT 1179.070 6.955 1179.350 7.325 ;
        RECT 1200.230 6.955 1200.510 7.325 ;
        RECT 1179.140 2.400 1179.280 6.955 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
      LAYER met3 ;
        RECT 1179.045 7.290 1179.375 7.305 ;
        RECT 1200.205 7.290 1200.535 7.305 ;
        RECT 1179.045 6.990 1200.535 7.290 ;
        RECT 1179.045 6.975 1179.375 6.990 ;
        RECT 1200.205 6.975 1200.535 6.990 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.090 14.010 1217.230 15.300 ;
        RECT 1216.860 13.870 1217.230 14.010 ;
        RECT 1216.860 10.725 1217.000 13.870 ;
        RECT 1196.550 10.355 1196.830 10.725 ;
        RECT 1216.790 10.355 1217.070 10.725 ;
        RECT 1196.620 2.400 1196.760 10.355 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
      LAYER met3 ;
        RECT 1196.525 10.690 1196.855 10.705 ;
        RECT 1216.765 10.690 1217.095 10.705 ;
        RECT 1196.525 10.390 1217.095 10.690 ;
        RECT 1196.525 10.375 1196.855 10.390 ;
        RECT 1216.765 10.375 1217.095 10.390 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.650 14.010 1233.790 15.300 ;
        RECT 1233.420 13.870 1233.790 14.010 ;
        RECT 1233.420 8.685 1233.560 13.870 ;
        RECT 1214.490 8.315 1214.770 8.685 ;
        RECT 1233.350 8.315 1233.630 8.685 ;
        RECT 1214.560 2.400 1214.700 8.315 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
      LAYER met3 ;
        RECT 1214.465 8.650 1214.795 8.665 ;
        RECT 1233.325 8.650 1233.655 8.665 ;
        RECT 1214.465 8.350 1233.655 8.650 ;
        RECT 1214.465 8.335 1214.795 8.350 ;
        RECT 1233.325 8.335 1233.655 8.350 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.210 14.010 1250.350 15.300 ;
        RECT 1249.980 13.870 1250.350 14.010 ;
        RECT 1249.980 12.085 1250.120 13.870 ;
        RECT 1231.970 11.715 1232.250 12.085 ;
        RECT 1249.910 11.715 1250.190 12.085 ;
        RECT 1232.040 2.400 1232.180 11.715 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
      LAYER met3 ;
        RECT 1231.945 12.050 1232.275 12.065 ;
        RECT 1249.885 12.050 1250.215 12.065 ;
        RECT 1231.945 11.750 1250.215 12.050 ;
        RECT 1231.945 11.735 1232.275 11.750 ;
        RECT 1249.885 11.735 1250.215 11.750 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.770 14.010 1266.910 15.300 ;
        RECT 1266.540 13.870 1266.910 14.010 ;
        RECT 1266.540 8.005 1266.680 13.870 ;
        RECT 1249.910 7.635 1250.190 8.005 ;
        RECT 1266.470 7.635 1266.750 8.005 ;
        RECT 1249.980 2.400 1250.120 7.635 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
      LAYER met3 ;
        RECT 1249.885 7.970 1250.215 7.985 ;
        RECT 1266.445 7.970 1266.775 7.985 ;
        RECT 1249.885 7.670 1266.775 7.970 ;
        RECT 1249.885 7.655 1250.215 7.670 ;
        RECT 1266.445 7.655 1266.775 7.670 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.330 14.010 1283.470 15.300 ;
        RECT 1283.100 13.870 1283.470 14.010 ;
        RECT 1283.100 8.005 1283.240 13.870 ;
        RECT 1267.390 7.635 1267.670 8.005 ;
        RECT 1283.030 7.635 1283.310 8.005 ;
        RECT 1267.460 2.400 1267.600 7.635 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
      LAYER met3 ;
        RECT 1267.365 7.970 1267.695 7.985 ;
        RECT 1283.005 7.970 1283.335 7.985 ;
        RECT 1267.365 7.670 1283.335 7.970 ;
        RECT 1267.365 7.655 1267.695 7.670 ;
        RECT 1283.005 7.655 1283.335 7.670 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.890 14.010 1300.030 15.300 ;
        RECT 1299.660 13.870 1300.030 14.010 ;
        RECT 1299.660 8.005 1299.800 13.870 ;
        RECT 1285.330 7.635 1285.610 8.005 ;
        RECT 1299.590 7.635 1299.870 8.005 ;
        RECT 1285.400 2.400 1285.540 7.635 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
      LAYER met3 ;
        RECT 1285.305 7.970 1285.635 7.985 ;
        RECT 1299.565 7.970 1299.895 7.985 ;
        RECT 1285.305 7.670 1299.895 7.970 ;
        RECT 1285.305 7.655 1285.635 7.670 ;
        RECT 1299.565 7.655 1299.895 7.670 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.450 14.010 1316.590 15.300 ;
        RECT 1316.220 13.870 1316.590 14.010 ;
        RECT 1316.220 8.005 1316.360 13.870 ;
        RECT 1303.270 7.635 1303.550 8.005 ;
        RECT 1316.150 7.635 1316.430 8.005 ;
        RECT 1303.340 2.400 1303.480 7.635 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
      LAYER met3 ;
        RECT 1303.245 7.970 1303.575 7.985 ;
        RECT 1316.125 7.970 1316.455 7.985 ;
        RECT 1303.245 7.670 1316.455 7.970 ;
        RECT 1303.245 7.655 1303.575 7.670 ;
        RECT 1316.125 7.655 1316.455 7.670 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.010 14.010 1333.150 15.300 ;
        RECT 1332.780 13.870 1333.150 14.010 ;
        RECT 1332.780 8.005 1332.920 13.870 ;
        RECT 1320.750 7.635 1321.030 8.005 ;
        RECT 1332.710 7.635 1332.990 8.005 ;
        RECT 1320.820 2.400 1320.960 7.635 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
      LAYER met3 ;
        RECT 1320.725 7.970 1321.055 7.985 ;
        RECT 1332.685 7.970 1333.015 7.985 ;
        RECT 1320.725 7.670 1333.015 7.970 ;
        RECT 1320.725 7.655 1321.055 7.670 ;
        RECT 1332.685 7.655 1333.015 7.670 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.850 14.010 736.990 15.300 ;
        RECT 736.620 13.870 736.990 14.010 ;
        RECT 736.620 3.925 736.760 13.870 ;
        RECT 682.270 3.555 682.550 3.925 ;
        RECT 736.550 3.555 736.830 3.925 ;
        RECT 682.340 2.400 682.480 3.555 ;
        RECT 682.130 -4.800 682.690 2.400 ;
      LAYER met3 ;
        RECT 682.245 3.890 682.575 3.905 ;
        RECT 736.525 3.890 736.855 3.905 ;
        RECT 682.245 3.590 736.855 3.890 ;
        RECT 682.245 3.575 682.575 3.590 ;
        RECT 736.525 3.575 736.855 3.590 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.570 14.010 1349.710 15.300 ;
        RECT 1349.340 13.870 1349.710 14.010 ;
        RECT 1349.340 6.645 1349.480 13.870 ;
        RECT 1338.690 6.275 1338.970 6.645 ;
        RECT 1349.270 6.275 1349.550 6.645 ;
        RECT 1338.760 2.400 1338.900 6.275 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
      LAYER met3 ;
        RECT 1338.665 6.610 1338.995 6.625 ;
        RECT 1349.245 6.610 1349.575 6.625 ;
        RECT 1338.665 6.310 1349.575 6.610 ;
        RECT 1338.665 6.295 1338.995 6.310 ;
        RECT 1349.245 6.295 1349.575 6.310 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.130 14.010 1366.270 15.300 ;
        RECT 1365.900 13.870 1366.270 14.010 ;
        RECT 1365.900 6.645 1366.040 13.870 ;
        RECT 1356.170 6.275 1356.450 6.645 ;
        RECT 1365.830 6.275 1366.110 6.645 ;
        RECT 1356.240 2.400 1356.380 6.275 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
      LAYER met3 ;
        RECT 1356.145 6.610 1356.475 6.625 ;
        RECT 1365.805 6.610 1366.135 6.625 ;
        RECT 1356.145 6.310 1366.135 6.610 ;
        RECT 1356.145 6.295 1356.475 6.310 ;
        RECT 1365.805 6.295 1366.135 6.310 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.690 14.010 1382.830 15.300 ;
        RECT 1382.460 13.870 1382.830 14.010 ;
        RECT 1382.460 5.965 1382.600 13.870 ;
        RECT 1374.110 5.595 1374.390 5.965 ;
        RECT 1382.390 5.595 1382.670 5.965 ;
        RECT 1374.180 2.400 1374.320 5.595 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
      LAYER met3 ;
        RECT 1374.085 5.930 1374.415 5.945 ;
        RECT 1382.365 5.930 1382.695 5.945 ;
        RECT 1374.085 5.630 1382.695 5.930 ;
        RECT 1374.085 5.615 1374.415 5.630 ;
        RECT 1382.365 5.615 1382.695 5.630 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.250 14.010 1399.390 15.300 ;
        RECT 1399.020 13.870 1399.390 14.010 ;
        RECT 1399.020 5.285 1399.160 13.870 ;
        RECT 1391.590 4.915 1391.870 5.285 ;
        RECT 1398.950 4.915 1399.230 5.285 ;
        RECT 1391.660 2.400 1391.800 4.915 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
      LAYER met3 ;
        RECT 1391.565 5.250 1391.895 5.265 ;
        RECT 1398.925 5.250 1399.255 5.265 ;
        RECT 1391.565 4.950 1399.255 5.250 ;
        RECT 1391.565 4.935 1391.895 4.950 ;
        RECT 1398.925 4.935 1399.255 4.950 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.810 14.690 1415.950 15.300 ;
        RECT 1415.810 14.550 1416.180 14.690 ;
        RECT 1416.040 6.645 1416.180 14.550 ;
        RECT 1409.530 6.275 1409.810 6.645 ;
        RECT 1415.970 6.275 1416.250 6.645 ;
        RECT 1409.600 2.400 1409.740 6.275 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
      LAYER met3 ;
        RECT 1409.505 6.610 1409.835 6.625 ;
        RECT 1415.945 6.610 1416.275 6.625 ;
        RECT 1409.505 6.310 1416.275 6.610 ;
        RECT 1409.505 6.295 1409.835 6.310 ;
        RECT 1415.945 6.295 1416.275 6.310 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.370 14.010 1432.510 15.300 ;
        RECT 1432.140 13.870 1432.510 14.010 ;
        RECT 1432.140 6.645 1432.280 13.870 ;
        RECT 1427.010 6.275 1427.290 6.645 ;
        RECT 1432.070 6.275 1432.350 6.645 ;
        RECT 1427.080 2.400 1427.220 6.275 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
      LAYER met3 ;
        RECT 1426.985 6.610 1427.315 6.625 ;
        RECT 1432.045 6.610 1432.375 6.625 ;
        RECT 1426.985 6.310 1432.375 6.610 ;
        RECT 1426.985 6.295 1427.315 6.310 ;
        RECT 1432.045 6.295 1432.375 6.310 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.930 14.010 1449.070 15.300 ;
        RECT 1447.320 13.870 1449.070 14.010 ;
        RECT 1444.810 1.770 1445.370 2.400 ;
        RECT 1447.320 1.770 1447.460 13.870 ;
        RECT 1444.810 1.630 1447.460 1.770 ;
        RECT 1444.810 -4.800 1445.370 1.630 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.490 14.010 1465.630 15.300 ;
        RECT 1462.960 13.870 1465.630 14.010 ;
        RECT 1462.960 2.400 1463.100 13.870 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.050 14.010 1482.190 15.300 ;
        RECT 1480.440 13.870 1482.190 14.010 ;
        RECT 1480.440 2.400 1480.580 13.870 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.610 14.010 1498.750 15.300 ;
        RECT 1498.380 13.870 1498.750 14.010 ;
        RECT 1498.380 2.400 1498.520 13.870 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.410 14.010 753.550 15.300 ;
        RECT 752.260 13.870 753.550 14.010 ;
        RECT 699.290 0.410 699.570 0.525 ;
        RECT 700.070 0.410 700.630 2.400 ;
        RECT 699.290 0.270 700.630 0.410 ;
        RECT 699.290 0.155 699.570 0.270 ;
        RECT 700.070 -4.800 700.630 0.270 ;
        RECT 751.730 0.410 752.010 0.525 ;
        RECT 752.260 0.410 752.400 13.870 ;
        RECT 751.730 0.270 752.400 0.410 ;
        RECT 751.730 0.155 752.010 0.270 ;
      LAYER met3 ;
        RECT 699.265 0.490 699.595 0.505 ;
        RECT 751.705 0.490 752.035 0.505 ;
        RECT 699.265 0.190 752.035 0.490 ;
        RECT 699.265 0.175 699.595 0.190 ;
        RECT 751.705 0.175 752.035 0.190 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.170 14.010 1515.310 15.300 ;
        RECT 1515.170 13.870 1516.000 14.010 ;
        RECT 1515.860 2.400 1516.000 13.870 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.730 14.010 1531.870 15.300 ;
        RECT 1531.730 13.870 1532.100 14.010 ;
        RECT 1531.960 1.770 1532.100 13.870 ;
        RECT 1533.590 1.770 1534.150 2.400 ;
        RECT 1531.960 1.630 1534.150 1.770 ;
        RECT 1533.590 -4.800 1534.150 1.630 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.290 14.010 1548.430 15.300 ;
        RECT 1548.290 13.870 1549.120 14.010 ;
        RECT 1548.980 1.770 1549.120 13.870 ;
        RECT 1551.070 1.770 1551.630 2.400 ;
        RECT 1548.980 1.630 1551.630 1.770 ;
        RECT 1551.070 -4.800 1551.630 1.630 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.850 14.010 1564.990 15.300 ;
        RECT 1564.850 13.870 1565.220 14.010 ;
        RECT 1565.080 6.645 1565.220 13.870 ;
        RECT 1565.010 6.275 1565.290 6.645 ;
        RECT 1569.150 6.275 1569.430 6.645 ;
        RECT 1569.220 2.400 1569.360 6.275 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
      LAYER met3 ;
        RECT 1564.985 6.610 1565.315 6.625 ;
        RECT 1569.125 6.610 1569.455 6.625 ;
        RECT 1564.985 6.310 1569.455 6.610 ;
        RECT 1564.985 6.295 1565.315 6.310 ;
        RECT 1569.125 6.295 1569.455 6.310 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.410 14.010 1581.550 15.300 ;
        RECT 1581.410 13.870 1586.840 14.010 ;
        RECT 1586.700 2.400 1586.840 13.870 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.970 14.010 1598.110 15.300 ;
        RECT 1597.970 13.870 1598.340 14.010 ;
        RECT 1598.200 6.645 1598.340 13.870 ;
        RECT 1598.130 6.275 1598.410 6.645 ;
        RECT 1604.570 6.275 1604.850 6.645 ;
        RECT 1604.640 2.400 1604.780 6.275 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
      LAYER met3 ;
        RECT 1598.105 6.610 1598.435 6.625 ;
        RECT 1604.545 6.610 1604.875 6.625 ;
        RECT 1598.105 6.310 1604.875 6.610 ;
        RECT 1598.105 6.295 1598.435 6.310 ;
        RECT 1604.545 6.295 1604.875 6.310 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.530 14.010 1614.670 15.300 ;
        RECT 1614.300 13.870 1614.670 14.010 ;
        RECT 1614.300 6.645 1614.440 13.870 ;
        RECT 1614.230 6.275 1614.510 6.645 ;
        RECT 1622.050 6.275 1622.330 6.645 ;
        RECT 1622.120 2.400 1622.260 6.275 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
      LAYER met3 ;
        RECT 1614.205 6.610 1614.535 6.625 ;
        RECT 1622.025 6.610 1622.355 6.625 ;
        RECT 1614.205 6.310 1622.355 6.610 ;
        RECT 1614.205 6.295 1614.535 6.310 ;
        RECT 1622.025 6.295 1622.355 6.310 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.090 14.010 1631.230 15.300 ;
        RECT 1631.090 13.870 1631.460 14.010 ;
        RECT 1631.320 5.965 1631.460 13.870 ;
        RECT 1631.250 5.595 1631.530 5.965 ;
        RECT 1639.990 5.595 1640.270 5.965 ;
        RECT 1640.060 2.400 1640.200 5.595 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
      LAYER met3 ;
        RECT 1631.225 5.930 1631.555 5.945 ;
        RECT 1639.965 5.930 1640.295 5.945 ;
        RECT 1631.225 5.630 1640.295 5.930 ;
        RECT 1631.225 5.615 1631.555 5.630 ;
        RECT 1639.965 5.615 1640.295 5.630 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.650 14.010 1647.790 15.300 ;
        RECT 1647.650 13.870 1648.020 14.010 ;
        RECT 1647.880 6.645 1648.020 13.870 ;
        RECT 1647.810 6.275 1648.090 6.645 ;
        RECT 1657.930 6.275 1658.210 6.645 ;
        RECT 1658.000 2.400 1658.140 6.275 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
      LAYER met3 ;
        RECT 1647.785 6.610 1648.115 6.625 ;
        RECT 1657.905 6.610 1658.235 6.625 ;
        RECT 1647.785 6.310 1658.235 6.610 ;
        RECT 1647.785 6.295 1648.115 6.310 ;
        RECT 1657.905 6.295 1658.235 6.310 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.210 14.010 1664.350 15.300 ;
        RECT 1664.210 13.870 1664.580 14.010 ;
        RECT 1664.440 5.965 1664.580 13.870 ;
        RECT 1664.370 5.595 1664.650 5.965 ;
        RECT 1675.410 5.595 1675.690 5.965 ;
        RECT 1675.480 2.400 1675.620 5.595 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
      LAYER met3 ;
        RECT 1664.345 5.930 1664.675 5.945 ;
        RECT 1675.385 5.930 1675.715 5.945 ;
        RECT 1664.345 5.630 1675.715 5.930 ;
        RECT 1664.345 5.615 1664.675 5.630 ;
        RECT 1675.385 5.615 1675.715 5.630 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.970 14.010 770.110 15.300 ;
        RECT 769.740 13.870 770.110 14.010 ;
        RECT 769.740 12.085 769.880 13.870 ;
        RECT 717.690 11.715 717.970 12.085 ;
        RECT 769.670 11.715 769.950 12.085 ;
        RECT 717.760 2.400 717.900 11.715 ;
        RECT 717.550 -4.800 718.110 2.400 ;
      LAYER met3 ;
        RECT 717.665 12.050 717.995 12.065 ;
        RECT 769.645 12.050 769.975 12.065 ;
        RECT 717.665 11.750 769.975 12.050 ;
        RECT 717.665 11.735 717.995 11.750 ;
        RECT 769.645 11.735 769.975 11.750 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.770 14.010 1680.910 15.300 ;
        RECT 1680.770 13.870 1681.140 14.010 ;
        RECT 1681.000 5.965 1681.140 13.870 ;
        RECT 1680.930 5.595 1681.210 5.965 ;
        RECT 1693.350 5.595 1693.630 5.965 ;
        RECT 1693.420 2.400 1693.560 5.595 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
      LAYER met3 ;
        RECT 1680.905 5.930 1681.235 5.945 ;
        RECT 1693.325 5.930 1693.655 5.945 ;
        RECT 1680.905 5.630 1693.655 5.930 ;
        RECT 1680.905 5.615 1681.235 5.630 ;
        RECT 1693.325 5.615 1693.655 5.630 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.330 14.010 1697.470 15.300 ;
        RECT 1697.100 13.870 1697.470 14.010 ;
        RECT 1697.100 5.965 1697.240 13.870 ;
        RECT 1697.030 5.595 1697.310 5.965 ;
        RECT 1710.830 5.595 1711.110 5.965 ;
        RECT 1710.900 2.400 1711.040 5.595 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
      LAYER met3 ;
        RECT 1697.005 5.930 1697.335 5.945 ;
        RECT 1710.805 5.930 1711.135 5.945 ;
        RECT 1697.005 5.630 1711.135 5.930 ;
        RECT 1697.005 5.615 1697.335 5.630 ;
        RECT 1710.805 5.615 1711.135 5.630 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.890 14.010 1714.030 15.300 ;
        RECT 1713.890 13.870 1714.260 14.010 ;
        RECT 1714.120 5.965 1714.260 13.870 ;
        RECT 1714.050 5.595 1714.330 5.965 ;
        RECT 1728.770 5.595 1729.050 5.965 ;
        RECT 1728.840 2.400 1728.980 5.595 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
      LAYER met3 ;
        RECT 1714.025 5.930 1714.355 5.945 ;
        RECT 1728.745 5.930 1729.075 5.945 ;
        RECT 1714.025 5.630 1729.075 5.930 ;
        RECT 1714.025 5.615 1714.355 5.630 ;
        RECT 1728.745 5.615 1729.075 5.630 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.450 14.125 1730.590 15.300 ;
        RECT 1730.380 13.755 1730.660 14.125 ;
        RECT 1746.250 13.755 1746.530 14.125 ;
        RECT 1746.320 2.400 1746.460 13.755 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
      LAYER met3 ;
        RECT 1730.355 14.090 1730.685 14.105 ;
        RECT 1746.225 14.090 1746.555 14.105 ;
        RECT 1730.355 13.790 1746.555 14.090 ;
        RECT 1730.355 13.775 1730.685 13.790 ;
        RECT 1746.225 13.775 1746.555 13.790 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.010 14.010 1747.150 15.300 ;
        RECT 1747.010 13.870 1747.380 14.010 ;
        RECT 1747.240 5.285 1747.380 13.870 ;
        RECT 1747.170 4.915 1747.450 5.285 ;
        RECT 1764.190 4.915 1764.470 5.285 ;
        RECT 1764.260 2.400 1764.400 4.915 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
      LAYER met3 ;
        RECT 1747.145 5.250 1747.475 5.265 ;
        RECT 1764.165 5.250 1764.495 5.265 ;
        RECT 1747.145 4.950 1764.495 5.250 ;
        RECT 1747.145 4.935 1747.475 4.950 ;
        RECT 1764.165 4.935 1764.495 4.950 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.570 14.125 1763.710 15.300 ;
        RECT 1763.500 13.755 1763.780 14.125 ;
        RECT 1781.670 13.755 1781.950 14.125 ;
        RECT 1781.740 2.400 1781.880 13.755 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
      LAYER met3 ;
        RECT 1763.475 14.090 1763.805 14.105 ;
        RECT 1781.645 14.090 1781.975 14.105 ;
        RECT 1763.475 13.790 1781.975 14.090 ;
        RECT 1763.475 13.775 1763.805 13.790 ;
        RECT 1781.645 13.775 1781.975 13.790 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.130 14.010 1780.270 15.300 ;
        RECT 1780.130 13.870 1780.500 14.010 ;
        RECT 1780.360 13.445 1780.500 13.870 ;
        RECT 1799.610 13.755 1799.890 14.125 ;
        RECT 1780.290 13.075 1780.570 13.445 ;
        RECT 1799.680 2.400 1799.820 13.755 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
      LAYER met3 ;
        RECT 1799.585 14.090 1799.915 14.105 ;
        RECT 1788.790 13.790 1799.915 14.090 ;
        RECT 1780.265 13.410 1780.595 13.425 ;
        RECT 1788.790 13.410 1789.090 13.790 ;
        RECT 1799.585 13.775 1799.915 13.790 ;
        RECT 1780.265 13.110 1789.090 13.410 ;
        RECT 1780.265 13.095 1780.595 13.110 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1796.600 14.520 1796.920 14.580 ;
        RECT 1816.610 14.520 1816.930 14.580 ;
        RECT 1796.600 14.380 1816.930 14.520 ;
        RECT 1796.600 14.320 1796.920 14.380 ;
        RECT 1816.610 14.320 1816.930 14.380 ;
      LAYER met2 ;
        RECT 1796.690 14.610 1796.830 15.300 ;
        RECT 1796.630 14.290 1796.890 14.610 ;
        RECT 1816.640 14.290 1816.900 14.610 ;
        RECT 1816.700 7.890 1816.840 14.290 ;
        RECT 1816.700 7.750 1817.760 7.890 ;
        RECT 1817.620 2.400 1817.760 7.750 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1813.390 7.720 1813.710 7.780 ;
        RECT 1834.090 7.720 1834.410 7.780 ;
        RECT 1813.390 7.580 1834.410 7.720 ;
        RECT 1813.390 7.520 1813.710 7.580 ;
        RECT 1834.090 7.520 1834.410 7.580 ;
      LAYER met2 ;
        RECT 1813.250 14.010 1813.390 15.300 ;
        RECT 1813.250 13.870 1813.620 14.010 ;
        RECT 1813.480 7.810 1813.620 13.870 ;
        RECT 1813.420 7.490 1813.680 7.810 ;
        RECT 1834.120 7.490 1834.380 7.810 ;
        RECT 1834.180 3.810 1834.320 7.490 ;
        RECT 1834.180 3.670 1835.240 3.810 ;
        RECT 1835.100 2.400 1835.240 3.670 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1829.720 14.520 1830.040 14.580 ;
        RECT 1850.190 14.520 1850.510 14.580 ;
        RECT 1829.720 14.380 1850.510 14.520 ;
        RECT 1829.720 14.320 1830.040 14.380 ;
        RECT 1850.190 14.320 1850.510 14.380 ;
      LAYER met2 ;
        RECT 1829.810 14.610 1829.950 15.300 ;
        RECT 1850.280 14.610 1850.880 14.690 ;
        RECT 1829.750 14.290 1830.010 14.610 ;
        RECT 1850.220 14.550 1850.880 14.610 ;
        RECT 1850.220 14.290 1850.480 14.550 ;
        RECT 1850.740 1.770 1850.880 14.550 ;
        RECT 1852.830 1.770 1853.390 2.400 ;
        RECT 1850.740 1.630 1853.390 1.770 ;
        RECT 1852.830 -4.800 1853.390 1.630 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.530 14.125 786.670 15.300 ;
        RECT 735.630 13.755 735.910 14.125 ;
        RECT 786.460 13.755 786.740 14.125 ;
        RECT 735.700 2.400 735.840 13.755 ;
        RECT 735.490 -4.800 736.050 2.400 ;
      LAYER met3 ;
        RECT 735.605 14.090 735.935 14.105 ;
        RECT 786.435 14.090 786.765 14.105 ;
        RECT 735.605 13.790 786.765 14.090 ;
        RECT 735.605 13.775 735.935 13.790 ;
        RECT 786.435 13.775 786.765 13.790 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1856.630 14.180 1856.950 14.240 ;
        RECT 1869.970 14.180 1870.290 14.240 ;
        RECT 1856.630 14.040 1870.290 14.180 ;
        RECT 1856.630 13.980 1856.950 14.040 ;
        RECT 1869.970 13.980 1870.290 14.040 ;
      LAYER met2 ;
        RECT 1846.370 14.125 1846.510 15.300 ;
        RECT 1856.660 14.125 1856.920 14.270 ;
        RECT 1846.300 13.755 1846.580 14.125 ;
        RECT 1856.650 13.755 1856.930 14.125 ;
        RECT 1870.000 13.950 1870.260 14.270 ;
        RECT 1870.060 7.210 1870.200 13.950 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.520 2.400 1870.660 7.070 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
      LAYER met3 ;
        RECT 1846.275 14.090 1846.605 14.105 ;
        RECT 1856.625 14.090 1856.955 14.105 ;
        RECT 1846.275 13.790 1856.955 14.090 ;
        RECT 1846.275 13.775 1846.605 13.790 ;
        RECT 1856.625 13.775 1856.955 13.790 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.930 14.690 1863.070 15.300 ;
        RECT 1862.700 14.550 1863.070 14.690 ;
        RECT 1862.700 14.125 1862.840 14.550 ;
        RECT 1862.630 13.755 1862.910 14.125 ;
        RECT 1887.470 12.650 1887.750 12.765 ;
        RECT 1887.470 12.510 1888.600 12.650 ;
        RECT 1887.470 12.395 1887.750 12.510 ;
        RECT 1888.460 2.400 1888.600 12.510 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
      LAYER met3 ;
        RECT 1887.190 15.450 1887.570 15.460 ;
        RECT 1863.310 15.150 1887.570 15.450 ;
        RECT 1862.605 14.090 1862.935 14.105 ;
        RECT 1863.310 14.090 1863.610 15.150 ;
        RECT 1887.190 15.140 1887.570 15.150 ;
        RECT 1862.605 13.790 1863.610 14.090 ;
        RECT 1862.605 13.775 1862.935 13.790 ;
        RECT 1887.445 12.740 1887.775 12.745 ;
        RECT 1887.190 12.730 1887.775 12.740 ;
        RECT 1887.190 12.430 1888.000 12.730 ;
        RECT 1887.190 12.420 1887.775 12.430 ;
        RECT 1887.445 12.415 1887.775 12.420 ;
      LAYER met4 ;
        RECT 1887.215 15.135 1887.545 15.465 ;
        RECT 1887.230 12.745 1887.530 15.135 ;
        RECT 1887.215 12.415 1887.545 12.745 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1879.400 14.180 1879.720 14.240 ;
        RECT 1904.470 14.180 1904.790 14.240 ;
        RECT 1879.400 14.040 1904.790 14.180 ;
        RECT 1879.400 13.980 1879.720 14.040 ;
        RECT 1904.470 13.980 1904.790 14.040 ;
      LAYER met2 ;
        RECT 1879.490 14.270 1879.630 15.300 ;
        RECT 1879.430 13.950 1879.690 14.270 ;
        RECT 1904.500 13.950 1904.760 14.270 ;
        RECT 1904.560 7.890 1904.700 13.950 ;
        RECT 1904.560 7.750 1906.080 7.890 ;
        RECT 1905.940 2.400 1906.080 7.750 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.050 14.125 1896.190 15.300 ;
        RECT 1895.980 13.755 1896.260 14.125 ;
        RECT 1923.810 13.755 1924.090 14.125 ;
        RECT 1923.880 2.400 1924.020 13.755 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
      LAYER met3 ;
        RECT 1895.955 14.090 1896.285 14.105 ;
        RECT 1923.785 14.090 1924.115 14.105 ;
        RECT 1895.955 13.790 1905.930 14.090 ;
        RECT 1895.955 13.775 1896.285 13.790 ;
        RECT 1905.630 13.410 1905.930 13.790 ;
        RECT 1920.350 13.790 1924.115 14.090 ;
        RECT 1920.350 13.410 1920.650 13.790 ;
        RECT 1923.785 13.775 1924.115 13.790 ;
        RECT 1905.630 13.110 1920.650 13.410 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.610 14.805 1912.750 15.300 ;
        RECT 1912.540 14.435 1912.820 14.805 ;
        RECT 1938.990 13.755 1939.270 14.125 ;
        RECT 1939.060 1.770 1939.200 13.755 ;
        RECT 1941.150 1.770 1941.710 2.400 ;
        RECT 1939.060 1.630 1941.710 1.770 ;
        RECT 1941.150 -4.800 1941.710 1.630 ;
      LAYER met3 ;
        RECT 1918.050 15.150 1939.050 15.450 ;
        RECT 1912.515 14.770 1912.845 14.785 ;
        RECT 1918.050 14.770 1918.350 15.150 ;
        RECT 1912.515 14.470 1918.350 14.770 ;
        RECT 1912.515 14.455 1912.845 14.470 ;
        RECT 1938.750 14.105 1939.050 15.150 ;
        RECT 1938.750 13.790 1939.295 14.105 ;
        RECT 1938.965 13.775 1939.295 13.790 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1929.080 14.520 1929.400 14.580 ;
        RECT 1959.210 14.520 1959.530 14.580 ;
        RECT 1929.080 14.380 1959.530 14.520 ;
        RECT 1929.080 14.320 1929.400 14.380 ;
        RECT 1959.210 14.320 1959.530 14.380 ;
      LAYER met2 ;
        RECT 1929.170 14.610 1929.310 15.300 ;
        RECT 1929.110 14.290 1929.370 14.610 ;
        RECT 1959.240 14.290 1959.500 14.610 ;
        RECT 1959.300 2.400 1959.440 14.290 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1945.640 14.180 1945.960 14.240 ;
        RECT 1967.490 14.180 1967.810 14.240 ;
        RECT 1945.640 14.040 1967.810 14.180 ;
        RECT 1945.640 13.980 1945.960 14.040 ;
        RECT 1967.490 13.980 1967.810 14.040 ;
      LAYER met2 ;
        RECT 1945.730 14.270 1945.870 15.300 ;
        RECT 1945.670 13.950 1945.930 14.270 ;
        RECT 1967.520 14.125 1967.780 14.270 ;
        RECT 1967.510 13.755 1967.790 14.125 ;
        RECT 1976.710 13.755 1976.990 14.125 ;
        RECT 1976.780 2.400 1976.920 13.755 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
      LAYER met3 ;
        RECT 1967.485 14.090 1967.815 14.105 ;
        RECT 1976.685 14.090 1977.015 14.105 ;
        RECT 1967.485 13.790 1977.015 14.090 ;
        RECT 1967.485 13.775 1967.815 13.790 ;
        RECT 1976.685 13.775 1977.015 13.790 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.290 14.805 1962.430 15.300 ;
        RECT 1962.220 14.435 1962.500 14.805 ;
        RECT 1994.190 13.330 1994.470 13.445 ;
        RECT 1994.190 13.190 1994.860 13.330 ;
        RECT 1994.190 13.075 1994.470 13.190 ;
        RECT 1994.720 2.400 1994.860 13.190 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
      LAYER met3 ;
        RECT 1962.195 14.770 1962.525 14.785 ;
        RECT 1962.195 14.470 1993.330 14.770 ;
        RECT 1962.195 14.455 1962.525 14.470 ;
        RECT 1993.030 13.410 1993.330 14.470 ;
        RECT 1994.165 13.410 1994.495 13.425 ;
        RECT 1993.030 13.110 1994.495 13.410 ;
        RECT 1994.165 13.095 1994.495 13.110 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1978.760 14.180 1979.080 14.240 ;
        RECT 2011.650 14.180 2011.970 14.240 ;
        RECT 1978.760 14.040 2011.970 14.180 ;
        RECT 1978.760 13.980 1979.080 14.040 ;
        RECT 2011.650 13.980 2011.970 14.040 ;
      LAYER met2 ;
        RECT 1978.850 14.270 1978.990 15.300 ;
        RECT 1978.790 13.950 1979.050 14.270 ;
        RECT 2011.680 13.950 2011.940 14.270 ;
        RECT 2011.740 7.890 2011.880 13.950 ;
        RECT 2011.740 7.750 2012.800 7.890 ;
        RECT 2012.660 2.400 2012.800 7.750 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.410 14.805 1995.550 15.300 ;
        RECT 1995.340 14.435 1995.620 14.805 ;
        RECT 2030.070 13.755 2030.350 14.125 ;
        RECT 2030.140 2.400 2030.280 13.755 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
      LAYER met3 ;
        RECT 2029.790 16.130 2030.170 16.140 ;
        RECT 2006.830 15.830 2030.170 16.130 ;
        RECT 1995.315 14.770 1995.645 14.785 ;
        RECT 2006.830 14.770 2007.130 15.830 ;
        RECT 2029.790 15.820 2030.170 15.830 ;
        RECT 1995.315 14.470 2007.130 14.770 ;
        RECT 1995.315 14.455 1995.645 14.470 ;
        RECT 2030.045 14.100 2030.375 14.105 ;
        RECT 2029.790 14.090 2030.375 14.100 ;
        RECT 2029.790 13.790 2030.600 14.090 ;
        RECT 2029.790 13.780 2030.375 13.790 ;
        RECT 2030.045 13.775 2030.375 13.780 ;
      LAYER met4 ;
        RECT 2029.815 15.815 2030.145 16.145 ;
        RECT 2029.830 14.105 2030.130 15.815 ;
        RECT 2029.815 13.775 2030.145 14.105 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.090 14.010 803.230 15.300 ;
        RECT 802.860 13.870 803.230 14.010 ;
        RECT 802.860 13.445 803.000 13.870 ;
        RECT 753.110 13.075 753.390 13.445 ;
        RECT 802.790 13.075 803.070 13.445 ;
        RECT 753.180 2.400 753.320 13.075 ;
        RECT 752.970 -4.800 753.530 2.400 ;
      LAYER met3 ;
        RECT 753.085 13.410 753.415 13.425 ;
        RECT 802.765 13.410 803.095 13.425 ;
        RECT 753.085 13.110 803.095 13.410 ;
        RECT 753.085 13.095 753.415 13.110 ;
        RECT 802.765 13.095 803.095 13.110 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2011.970 14.805 2012.110 15.300 ;
        RECT 2011.900 14.435 2012.180 14.805 ;
        RECT 2048.010 13.755 2048.290 14.125 ;
        RECT 2048.080 2.400 2048.220 13.755 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
      LAYER met3 ;
        RECT 2014.650 15.150 2043.930 15.450 ;
        RECT 2011.875 14.770 2012.205 14.785 ;
        RECT 2014.650 14.770 2014.950 15.150 ;
        RECT 2011.875 14.470 2014.950 14.770 ;
        RECT 2011.875 14.455 2012.205 14.470 ;
        RECT 2043.630 14.090 2043.930 15.150 ;
        RECT 2047.985 14.090 2048.315 14.105 ;
        RECT 2043.630 13.790 2048.315 14.090 ;
        RECT 2047.985 13.775 2048.315 13.790 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.530 14.010 2028.670 15.300 ;
        RECT 2028.300 13.870 2028.670 14.010 ;
        RECT 2028.300 1.885 2028.440 13.870 ;
        RECT 2028.230 1.515 2028.510 1.885 ;
        RECT 2064.110 1.770 2064.390 1.885 ;
        RECT 2065.350 1.770 2065.910 2.400 ;
        RECT 2064.110 1.630 2065.910 1.770 ;
        RECT 2064.110 1.515 2064.390 1.630 ;
        RECT 2065.350 -4.800 2065.910 1.630 ;
      LAYER met3 ;
        RECT 2028.205 1.850 2028.535 1.865 ;
        RECT 2064.085 1.850 2064.415 1.865 ;
        RECT 2028.205 1.550 2064.415 1.850 ;
        RECT 2028.205 1.535 2028.535 1.550 ;
        RECT 2064.085 1.535 2064.415 1.550 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.090 14.805 2045.230 15.300 ;
        RECT 2045.020 14.435 2045.300 14.805 ;
        RECT 2082.970 13.755 2083.250 14.125 ;
        RECT 2083.040 5.170 2083.180 13.755 ;
        RECT 2083.040 5.030 2083.640 5.170 ;
        RECT 2083.500 2.400 2083.640 5.030 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
      LAYER met3 ;
        RECT 2044.995 14.770 2045.325 14.785 ;
        RECT 2044.995 14.470 2074.290 14.770 ;
        RECT 2044.995 14.455 2045.325 14.470 ;
        RECT 2073.990 14.090 2074.290 14.470 ;
        RECT 2082.945 14.090 2083.275 14.105 ;
        RECT 2073.990 13.790 2083.275 14.090 ;
        RECT 2082.945 13.775 2083.275 13.790 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.650 14.010 2061.790 15.300 ;
        RECT 2061.650 13.870 2062.020 14.010 ;
        RECT 2061.880 4.605 2062.020 13.870 ;
        RECT 2061.810 4.235 2062.090 4.605 ;
        RECT 2100.910 4.235 2101.190 4.605 ;
        RECT 2100.980 2.400 2101.120 4.235 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
      LAYER met3 ;
        RECT 2061.785 4.570 2062.115 4.585 ;
        RECT 2100.885 4.570 2101.215 4.585 ;
        RECT 2061.785 4.270 2101.215 4.570 ;
        RECT 2061.785 4.255 2062.115 4.270 ;
        RECT 2100.885 4.255 2101.215 4.270 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.210 14.010 2078.350 15.300 ;
        RECT 2078.210 13.870 2078.580 14.010 ;
        RECT 2078.440 6.645 2078.580 13.870 ;
        RECT 2078.370 6.275 2078.650 6.645 ;
        RECT 2118.850 6.275 2119.130 6.645 ;
        RECT 2118.920 2.400 2119.060 6.275 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
      LAYER met3 ;
        RECT 2078.345 6.610 2078.675 6.625 ;
        RECT 2118.825 6.610 2119.155 6.625 ;
        RECT 2078.345 6.310 2119.155 6.610 ;
        RECT 2078.345 6.295 2078.675 6.310 ;
        RECT 2118.825 6.295 2119.155 6.310 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.770 14.010 2094.910 15.300 ;
        RECT 2094.770 13.870 2095.140 14.010 ;
        RECT 2095.000 10.045 2095.140 13.870 ;
        RECT 2094.930 9.675 2095.210 10.045 ;
        RECT 2136.330 9.675 2136.610 10.045 ;
        RECT 2136.400 2.400 2136.540 9.675 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
      LAYER met3 ;
        RECT 2094.905 10.010 2095.235 10.025 ;
        RECT 2136.305 10.010 2136.635 10.025 ;
        RECT 2094.905 9.710 2136.635 10.010 ;
        RECT 2094.905 9.695 2095.235 9.710 ;
        RECT 2136.305 9.695 2136.635 9.710 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2111.010 0.580 2111.330 0.640 ;
        RECT 2155.170 0.580 2155.490 0.640 ;
        RECT 2111.010 0.440 2155.490 0.580 ;
        RECT 2111.010 0.380 2111.330 0.440 ;
        RECT 2155.170 0.380 2155.490 0.440 ;
      LAYER met2 ;
        RECT 2111.330 14.010 2111.470 15.300 ;
        RECT 2111.100 13.870 2111.470 14.010 ;
        RECT 2111.100 0.670 2111.240 13.870 ;
        RECT 2111.040 0.350 2111.300 0.670 ;
        RECT 2154.130 0.410 2154.690 2.400 ;
        RECT 2155.200 0.410 2155.460 0.670 ;
        RECT 2154.130 0.350 2155.460 0.410 ;
        RECT 2154.130 0.270 2155.400 0.350 ;
        RECT 2154.130 -4.800 2154.690 0.270 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.890 14.010 2128.030 15.300 ;
        RECT 2127.890 13.870 2128.260 14.010 ;
        RECT 2128.120 6.645 2128.260 13.870 ;
        RECT 2128.050 6.275 2128.330 6.645 ;
        RECT 2172.210 6.275 2172.490 6.645 ;
        RECT 2172.280 2.400 2172.420 6.275 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
      LAYER met3 ;
        RECT 2128.025 6.610 2128.355 6.625 ;
        RECT 2172.185 6.610 2172.515 6.625 ;
        RECT 2128.025 6.310 2172.515 6.610 ;
        RECT 2128.025 6.295 2128.355 6.310 ;
        RECT 2172.185 6.295 2172.515 6.310 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.450 14.010 2144.590 15.300 ;
        RECT 2144.450 13.870 2144.820 14.010 ;
        RECT 2144.680 1.885 2144.820 13.870 ;
        RECT 2144.610 1.515 2144.890 1.885 ;
        RECT 2187.390 1.770 2187.670 1.885 ;
        RECT 2189.550 1.770 2190.110 2.400 ;
        RECT 2187.390 1.630 2190.110 1.770 ;
        RECT 2187.390 1.515 2187.670 1.630 ;
        RECT 2189.550 -4.800 2190.110 1.630 ;
      LAYER met3 ;
        RECT 2144.585 1.850 2144.915 1.865 ;
        RECT 2187.365 1.850 2187.695 1.865 ;
        RECT 2144.585 1.550 2187.695 1.850 ;
        RECT 2144.585 1.535 2144.915 1.550 ;
        RECT 2187.365 1.535 2187.695 1.550 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.010 14.010 2161.150 15.300 ;
        RECT 2161.010 13.870 2161.380 14.010 ;
        RECT 2161.240 5.965 2161.380 13.870 ;
        RECT 2161.170 5.595 2161.450 5.965 ;
        RECT 2207.630 5.595 2207.910 5.965 ;
        RECT 2207.700 2.400 2207.840 5.595 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
      LAYER met3 ;
        RECT 2161.145 5.930 2161.475 5.945 ;
        RECT 2207.605 5.930 2207.935 5.945 ;
        RECT 2161.145 5.630 2207.935 5.930 ;
        RECT 2161.145 5.615 2161.475 5.630 ;
        RECT 2207.605 5.615 2207.935 5.630 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.650 14.010 819.790 15.300 ;
        RECT 819.420 13.870 819.790 14.010 ;
        RECT 819.420 10.725 819.560 13.870 ;
        RECT 771.050 10.355 771.330 10.725 ;
        RECT 819.350 10.355 819.630 10.725 ;
        RECT 771.120 2.400 771.260 10.355 ;
        RECT 770.910 -4.800 771.470 2.400 ;
      LAYER met3 ;
        RECT 771.025 10.690 771.355 10.705 ;
        RECT 819.325 10.690 819.655 10.705 ;
        RECT 771.025 10.390 819.655 10.690 ;
        RECT 771.025 10.375 771.355 10.390 ;
        RECT 819.325 10.375 819.655 10.390 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.570 14.010 2177.710 15.300 ;
        RECT 2177.570 13.870 2177.940 14.010 ;
        RECT 2177.800 11.405 2177.940 13.870 ;
        RECT 2177.730 11.035 2178.010 11.405 ;
        RECT 2225.110 11.035 2225.390 11.405 ;
        RECT 2225.180 2.400 2225.320 11.035 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
      LAYER met3 ;
        RECT 2177.705 11.370 2178.035 11.385 ;
        RECT 2225.085 11.370 2225.415 11.385 ;
        RECT 2177.705 11.070 2225.415 11.370 ;
        RECT 2177.705 11.055 2178.035 11.070 ;
        RECT 2225.085 11.055 2225.415 11.070 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2193.810 0.920 2194.130 0.980 ;
        RECT 2242.110 0.920 2242.430 0.980 ;
        RECT 2193.810 0.780 2242.430 0.920 ;
        RECT 2193.810 0.720 2194.130 0.780 ;
        RECT 2242.110 0.720 2242.430 0.780 ;
      LAYER met2 ;
        RECT 2194.130 14.010 2194.270 15.300 ;
        RECT 2193.900 13.870 2194.270 14.010 ;
        RECT 2193.900 1.010 2194.040 13.870 ;
        RECT 2242.910 1.090 2243.470 2.400 ;
        RECT 2242.200 1.010 2243.470 1.090 ;
        RECT 2193.840 0.690 2194.100 1.010 ;
        RECT 2242.140 0.950 2243.470 1.010 ;
        RECT 2242.140 0.690 2242.400 0.950 ;
        RECT 2242.910 -4.800 2243.470 0.950 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.690 14.010 2210.830 15.300 ;
        RECT 2210.690 13.870 2211.060 14.010 ;
        RECT 2210.920 12.765 2211.060 13.870 ;
        RECT 2210.850 12.395 2211.130 12.765 ;
        RECT 2260.530 12.395 2260.810 12.765 ;
        RECT 2260.600 2.400 2260.740 12.395 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
      LAYER met3 ;
        RECT 2210.825 12.730 2211.155 12.745 ;
        RECT 2260.505 12.730 2260.835 12.745 ;
        RECT 2210.825 12.430 2260.835 12.730 ;
        RECT 2210.825 12.415 2211.155 12.430 ;
        RECT 2260.505 12.415 2260.835 12.430 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2227.250 14.010 2227.390 15.300 ;
        RECT 2227.250 13.870 2227.620 14.010 ;
        RECT 2227.480 11.405 2227.620 13.870 ;
        RECT 2227.410 11.035 2227.690 11.405 ;
        RECT 2278.470 11.035 2278.750 11.405 ;
        RECT 2278.540 2.400 2278.680 11.035 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
      LAYER met3 ;
        RECT 2227.385 11.370 2227.715 11.385 ;
        RECT 2278.445 11.370 2278.775 11.385 ;
        RECT 2227.385 11.070 2278.775 11.370 ;
        RECT 2227.385 11.055 2227.715 11.070 ;
        RECT 2278.445 11.055 2278.775 11.070 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.810 14.010 2243.950 15.300 ;
        RECT 2243.810 13.870 2244.180 14.010 ;
        RECT 2244.040 10.045 2244.180 13.870 ;
        RECT 2243.970 9.675 2244.250 10.045 ;
        RECT 2295.950 9.675 2296.230 10.045 ;
        RECT 2296.020 2.400 2296.160 9.675 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
      LAYER met3 ;
        RECT 2243.945 10.010 2244.275 10.025 ;
        RECT 2295.925 10.010 2296.255 10.025 ;
        RECT 2243.945 9.710 2296.255 10.010 ;
        RECT 2243.945 9.695 2244.275 9.710 ;
        RECT 2295.925 9.695 2296.255 9.710 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.370 14.805 2260.510 15.300 ;
        RECT 2260.300 14.435 2260.580 14.805 ;
        RECT 2313.430 13.330 2313.710 13.445 ;
        RECT 2313.430 13.190 2314.100 13.330 ;
        RECT 2313.430 13.075 2313.710 13.190 ;
        RECT 2313.960 2.400 2314.100 13.190 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
      LAYER met3 ;
        RECT 2313.150 18.170 2313.530 18.180 ;
        RECT 2264.430 17.870 2313.530 18.170 ;
        RECT 2260.275 14.770 2260.605 14.785 ;
        RECT 2264.430 14.770 2264.730 17.870 ;
        RECT 2313.150 17.860 2313.530 17.870 ;
        RECT 2260.275 14.470 2264.730 14.770 ;
        RECT 2260.275 14.455 2260.605 14.470 ;
        RECT 2313.405 13.420 2313.735 13.425 ;
        RECT 2313.150 13.410 2313.735 13.420 ;
        RECT 2313.150 13.110 2313.960 13.410 ;
        RECT 2313.150 13.100 2313.735 13.110 ;
        RECT 2313.405 13.095 2313.735 13.100 ;
      LAYER met4 ;
        RECT 2313.175 17.855 2313.505 18.185 ;
        RECT 2313.190 13.425 2313.490 17.855 ;
        RECT 2313.175 13.095 2313.505 13.425 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.930 14.805 2277.070 15.300 ;
        RECT 2276.860 14.435 2277.140 14.805 ;
        RECT 2331.370 12.395 2331.650 12.765 ;
        RECT 2331.440 2.400 2331.580 12.395 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
      LAYER met3 ;
        RECT 2331.550 16.130 2331.930 16.140 ;
        RECT 2276.850 15.830 2331.930 16.130 ;
        RECT 2276.850 14.785 2277.150 15.830 ;
        RECT 2331.550 15.820 2331.930 15.830 ;
        RECT 2276.835 14.455 2277.165 14.785 ;
        RECT 2331.345 12.740 2331.675 12.745 ;
        RECT 2331.345 12.730 2331.930 12.740 ;
        RECT 2331.120 12.430 2331.930 12.730 ;
        RECT 2331.345 12.420 2331.930 12.430 ;
        RECT 2331.345 12.415 2331.675 12.420 ;
      LAYER met4 ;
        RECT 2331.575 15.815 2331.905 16.145 ;
        RECT 2331.590 12.745 2331.890 15.815 ;
        RECT 2331.575 12.415 2331.905 12.745 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2293.490 14.805 2293.630 15.300 ;
        RECT 2293.420 14.435 2293.700 14.805 ;
        RECT 2349.310 13.755 2349.590 14.125 ;
        RECT 2349.380 2.400 2349.520 13.755 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
      LAYER met3 ;
        RECT 2293.395 14.770 2293.725 14.785 ;
        RECT 2293.395 14.470 2297.850 14.770 ;
        RECT 2293.395 14.455 2293.725 14.470 ;
        RECT 2297.550 14.090 2297.850 14.470 ;
        RECT 2349.285 14.090 2349.615 14.105 ;
        RECT 2297.550 13.790 2318.090 14.090 ;
        RECT 2317.790 13.410 2318.090 13.790 ;
        RECT 2321.470 13.790 2349.615 14.090 ;
        RECT 2321.470 13.410 2321.770 13.790 ;
        RECT 2349.285 13.775 2349.615 13.790 ;
        RECT 2317.790 13.110 2321.770 13.410 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2310.190 6.700 2310.510 6.760 ;
        RECT 2310.190 6.560 2331.580 6.700 ;
        RECT 2310.190 6.500 2310.510 6.560 ;
        RECT 2331.440 6.360 2331.580 6.560 ;
        RECT 2366.770 6.360 2367.090 6.420 ;
        RECT 2331.440 6.220 2367.090 6.360 ;
        RECT 2366.770 6.160 2367.090 6.220 ;
      LAYER met2 ;
        RECT 2310.050 13.870 2310.190 15.300 ;
        RECT 2310.050 13.730 2310.420 13.870 ;
        RECT 2310.280 6.790 2310.420 13.730 ;
        RECT 2310.220 6.470 2310.480 6.790 ;
        RECT 2366.800 6.130 2367.060 6.450 ;
        RECT 2366.860 3.130 2367.000 6.130 ;
        RECT 2366.860 2.990 2367.460 3.130 ;
        RECT 2367.320 2.400 2367.460 2.990 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2326.610 13.870 2326.750 15.300 ;
        RECT 2326.610 13.730 2326.980 13.870 ;
        RECT 2326.840 2.565 2326.980 13.730 ;
        RECT 2326.770 2.195 2327.050 2.565 ;
        RECT 2381.970 2.450 2382.250 2.565 ;
        RECT 2381.970 2.310 2382.640 2.450 ;
        RECT 2381.970 2.195 2382.250 2.310 ;
        RECT 2382.500 1.770 2382.640 2.310 ;
        RECT 2384.590 1.770 2385.150 2.400 ;
        RECT 2382.500 1.630 2385.150 1.770 ;
        RECT 2384.590 -4.800 2385.150 1.630 ;
      LAYER met3 ;
        RECT 2326.745 2.530 2327.075 2.545 ;
        RECT 2381.945 2.530 2382.275 2.545 ;
        RECT 2326.745 2.230 2382.275 2.530 ;
        RECT 2326.745 2.215 2327.075 2.230 ;
        RECT 2381.945 2.215 2382.275 2.230 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.210 14.010 836.350 15.300 ;
        RECT 835.980 13.870 836.350 14.010 ;
        RECT 835.980 8.685 836.120 13.870 ;
        RECT 788.990 8.315 789.270 8.685 ;
        RECT 835.910 8.315 836.190 8.685 ;
        RECT 789.060 2.400 789.200 8.315 ;
        RECT 788.850 -4.800 789.410 2.400 ;
      LAYER met3 ;
        RECT 788.965 8.650 789.295 8.665 ;
        RECT 835.885 8.650 836.215 8.665 ;
        RECT 788.965 8.350 836.215 8.650 ;
        RECT 788.965 8.335 789.295 8.350 ;
        RECT 835.885 8.335 836.215 8.350 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.690 14.010 692.830 15.300 ;
        RECT 692.460 13.870 692.830 14.010 ;
        RECT 634.960 2.990 636.020 3.130 ;
        RECT 634.960 2.400 635.100 2.990 ;
        RECT 634.750 -4.800 635.310 2.400 ;
        RECT 635.880 1.885 636.020 2.990 ;
        RECT 692.460 1.885 692.600 13.870 ;
        RECT 635.810 1.515 636.090 1.885 ;
        RECT 692.390 1.515 692.670 1.885 ;
      LAYER met3 ;
        RECT 635.785 1.850 636.115 1.865 ;
        RECT 692.365 1.850 692.695 1.865 ;
        RECT 635.785 1.550 692.695 1.850 ;
        RECT 635.785 1.535 636.115 1.550 ;
        RECT 692.365 1.535 692.695 1.550 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2348.690 14.010 2348.830 15.300 ;
        RECT 2348.690 13.870 2349.060 14.010 ;
        RECT 2348.920 10.045 2349.060 13.870 ;
        RECT 2348.850 9.675 2349.130 10.045 ;
        RECT 2408.650 9.675 2408.930 10.045 ;
        RECT 2408.720 2.400 2408.860 9.675 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
      LAYER met3 ;
        RECT 2348.825 10.010 2349.155 10.025 ;
        RECT 2408.625 10.010 2408.955 10.025 ;
        RECT 2348.825 9.710 2408.955 10.010 ;
        RECT 2348.825 9.695 2349.155 9.710 ;
        RECT 2408.625 9.695 2408.955 9.710 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2394.370 14.180 2394.690 14.240 ;
        RECT 2426.110 14.180 2426.430 14.240 ;
        RECT 2394.370 14.040 2426.430 14.180 ;
        RECT 2394.370 13.980 2394.690 14.040 ;
        RECT 2426.110 13.980 2426.430 14.040 ;
        RECT 2365.390 6.700 2365.710 6.760 ;
        RECT 2394.370 6.700 2394.690 6.760 ;
        RECT 2365.390 6.560 2394.690 6.700 ;
        RECT 2365.390 6.500 2365.710 6.560 ;
        RECT 2394.370 6.500 2394.690 6.560 ;
      LAYER met2 ;
        RECT 2365.250 14.010 2365.390 15.300 ;
        RECT 2365.250 13.870 2365.620 14.010 ;
        RECT 2394.400 13.950 2394.660 14.270 ;
        RECT 2426.140 13.950 2426.400 14.270 ;
        RECT 2365.480 6.790 2365.620 13.870 ;
        RECT 2394.460 6.790 2394.600 13.950 ;
        RECT 2365.420 6.470 2365.680 6.790 ;
        RECT 2394.400 6.470 2394.660 6.790 ;
        RECT 2426.200 2.400 2426.340 13.950 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.810 14.010 2381.950 15.300 ;
        RECT 2381.580 13.870 2381.950 14.010 ;
        RECT 2381.580 0.525 2381.720 13.870 ;
        RECT 2381.510 0.155 2381.790 0.525 ;
        RECT 2443.930 0.410 2444.490 2.400 ;
        RECT 2444.990 0.410 2445.270 0.525 ;
        RECT 2443.930 0.270 2445.270 0.410 ;
        RECT 2443.930 -4.800 2444.490 0.270 ;
        RECT 2444.990 0.155 2445.270 0.270 ;
      LAYER met3 ;
        RECT 2381.485 0.490 2381.815 0.505 ;
        RECT 2444.965 0.490 2445.295 0.505 ;
        RECT 2381.485 0.190 2445.295 0.490 ;
        RECT 2381.485 0.175 2381.815 0.190 ;
        RECT 2444.965 0.175 2445.295 0.190 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2398.510 6.700 2398.830 6.760 ;
        RECT 2460.150 6.700 2460.470 6.760 ;
        RECT 2398.510 6.560 2460.470 6.700 ;
        RECT 2398.510 6.500 2398.830 6.560 ;
        RECT 2460.150 6.500 2460.470 6.560 ;
      LAYER met2 ;
        RECT 2398.370 14.010 2398.510 15.300 ;
        RECT 2398.370 13.870 2398.740 14.010 ;
        RECT 2398.600 6.790 2398.740 13.870 ;
        RECT 2398.540 6.470 2398.800 6.790 ;
        RECT 2460.180 6.470 2460.440 6.790 ;
        RECT 2460.240 3.810 2460.380 6.470 ;
        RECT 2460.240 3.670 2461.760 3.810 ;
        RECT 2461.620 2.400 2461.760 3.670 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2414.610 3.300 2414.930 3.360 ;
        RECT 2479.470 3.300 2479.790 3.360 ;
        RECT 2414.610 3.160 2479.790 3.300 ;
        RECT 2414.610 3.100 2414.930 3.160 ;
        RECT 2479.470 3.100 2479.790 3.160 ;
      LAYER met2 ;
        RECT 2414.930 14.010 2415.070 15.300 ;
        RECT 2414.700 13.870 2415.070 14.010 ;
        RECT 2414.700 3.390 2414.840 13.870 ;
        RECT 2414.640 3.070 2414.900 3.390 ;
        RECT 2479.500 3.070 2479.760 3.390 ;
        RECT 2479.560 2.400 2479.700 3.070 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.490 14.010 2431.630 15.300 ;
        RECT 2430.800 13.870 2431.630 14.010 ;
        RECT 2430.800 1.885 2430.940 13.870 ;
        RECT 2430.730 1.515 2431.010 1.885 ;
        RECT 2494.670 1.770 2494.950 1.885 ;
        RECT 2496.830 1.770 2497.390 2.400 ;
        RECT 2494.670 1.630 2497.390 1.770 ;
        RECT 2494.670 1.515 2494.950 1.630 ;
        RECT 2496.830 -4.800 2497.390 1.630 ;
      LAYER met3 ;
        RECT 2430.705 1.850 2431.035 1.865 ;
        RECT 2494.645 1.850 2494.975 1.865 ;
        RECT 2430.705 1.550 2494.975 1.850 ;
        RECT 2430.705 1.535 2431.035 1.550 ;
        RECT 2494.645 1.535 2494.975 1.550 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2448.050 14.010 2448.190 15.300 ;
        RECT 2448.050 13.870 2448.420 14.010 ;
        RECT 2448.280 0.525 2448.420 13.870 ;
        RECT 2448.210 0.155 2448.490 0.525 ;
        RECT 2514.770 0.410 2515.330 2.400 ;
        RECT 2515.830 0.410 2516.110 0.525 ;
        RECT 2514.770 0.270 2516.110 0.410 ;
        RECT 2514.770 -4.800 2515.330 0.270 ;
        RECT 2515.830 0.155 2516.110 0.270 ;
      LAYER met3 ;
        RECT 2448.185 0.490 2448.515 0.505 ;
        RECT 2515.805 0.490 2516.135 0.505 ;
        RECT 2448.185 0.190 2516.135 0.490 ;
        RECT 2448.185 0.175 2448.515 0.190 ;
        RECT 2515.805 0.175 2516.135 0.190 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.610 14.010 2464.750 15.300 ;
        RECT 2464.610 13.870 2464.980 14.010 ;
        RECT 2464.840 2.565 2464.980 13.870 ;
        RECT 2464.770 2.195 2465.050 2.565 ;
        RECT 2532.250 1.770 2532.810 2.400 ;
        RECT 2533.310 2.195 2533.590 2.565 ;
        RECT 2533.380 1.770 2533.520 2.195 ;
        RECT 2532.250 1.630 2533.520 1.770 ;
        RECT 2532.250 -4.800 2532.810 1.630 ;
      LAYER met3 ;
        RECT 2464.745 2.530 2465.075 2.545 ;
        RECT 2533.285 2.530 2533.615 2.545 ;
        RECT 2464.745 2.230 2533.615 2.530 ;
        RECT 2464.745 2.215 2465.075 2.230 ;
        RECT 2533.285 2.215 2533.615 2.230 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2481.310 6.700 2481.630 6.760 ;
        RECT 2548.010 6.700 2548.330 6.760 ;
        RECT 2481.310 6.560 2548.330 6.700 ;
        RECT 2481.310 6.500 2481.630 6.560 ;
        RECT 2548.010 6.500 2548.330 6.560 ;
      LAYER met2 ;
        RECT 2481.170 14.010 2481.310 15.300 ;
        RECT 2481.170 13.870 2481.540 14.010 ;
        RECT 2481.400 6.790 2481.540 13.870 ;
        RECT 2481.340 6.470 2481.600 6.790 ;
        RECT 2548.040 6.470 2548.300 6.790 ;
        RECT 2548.100 1.770 2548.240 6.470 ;
        RECT 2550.190 1.770 2550.750 2.400 ;
        RECT 2548.100 1.630 2550.750 1.770 ;
        RECT 2550.190 -4.800 2550.750 1.630 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2497.410 3.300 2497.730 3.360 ;
        RECT 2497.410 3.100 2497.870 3.300 ;
        RECT 2497.730 1.600 2497.870 3.100 ;
        RECT 2566.870 1.600 2567.190 1.660 ;
        RECT 2497.730 1.460 2567.190 1.600 ;
        RECT 2566.870 1.400 2567.190 1.460 ;
      LAYER met2 ;
        RECT 2497.730 14.010 2497.870 15.300 ;
        RECT 2497.500 13.870 2497.870 14.010 ;
        RECT 2497.500 3.390 2497.640 13.870 ;
        RECT 2497.440 3.070 2497.700 3.390 ;
        RECT 2567.670 1.770 2568.230 2.400 ;
        RECT 2566.960 1.690 2568.230 1.770 ;
        RECT 2566.900 1.630 2568.230 1.690 ;
        RECT 2566.900 1.370 2567.160 1.630 ;
        RECT 2567.670 -4.800 2568.230 1.630 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.290 14.010 858.430 15.300 ;
        RECT 858.060 13.870 858.430 14.010 ;
        RECT 858.060 12.765 858.200 13.870 ;
        RECT 812.450 12.395 812.730 12.765 ;
        RECT 857.990 12.395 858.270 12.765 ;
        RECT 812.520 2.400 812.660 12.395 ;
        RECT 812.310 -4.800 812.870 2.400 ;
      LAYER met3 ;
        RECT 812.425 12.730 812.755 12.745 ;
        RECT 857.965 12.730 858.295 12.745 ;
        RECT 812.425 12.430 858.295 12.730 ;
        RECT 812.425 12.415 812.755 12.430 ;
        RECT 857.965 12.415 858.295 12.430 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.290 14.010 2514.430 15.300 ;
        RECT 2513.600 13.870 2514.430 14.010 ;
        RECT 2513.600 1.205 2513.740 13.870 ;
        RECT 2585.750 2.875 2586.030 3.245 ;
        RECT 2585.820 2.400 2585.960 2.875 ;
        RECT 2513.530 0.835 2513.810 1.205 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
      LAYER met3 ;
        RECT 2585.725 3.210 2586.055 3.225 ;
        RECT 2578.150 2.910 2586.055 3.210 ;
        RECT 2513.505 1.170 2513.835 1.185 ;
        RECT 2578.150 1.170 2578.450 2.910 ;
        RECT 2585.725 2.895 2586.055 2.910 ;
        RECT 2513.505 0.870 2578.450 1.170 ;
        RECT 2513.505 0.855 2513.835 0.870 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2603.670 3.300 2603.990 3.360 ;
        RECT 2594.330 3.160 2603.990 3.300 ;
        RECT 2530.990 1.940 2531.310 2.000 ;
        RECT 2594.330 1.940 2594.470 3.160 ;
        RECT 2603.670 3.100 2603.990 3.160 ;
        RECT 2530.990 1.800 2594.470 1.940 ;
        RECT 2530.990 1.740 2531.310 1.800 ;
      LAYER met2 ;
        RECT 2530.850 14.010 2530.990 15.300 ;
        RECT 2530.850 13.870 2531.220 14.010 ;
        RECT 2531.080 2.030 2531.220 13.870 ;
        RECT 2603.700 3.070 2603.960 3.390 ;
        RECT 2603.760 2.400 2603.900 3.070 ;
        RECT 2531.020 1.710 2531.280 2.030 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.410 14.125 2547.550 15.300 ;
        RECT 2547.340 13.755 2547.620 14.125 ;
        RECT 2621.170 13.755 2621.450 14.125 ;
        RECT 2621.240 2.400 2621.380 13.755 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
      LAYER met3 ;
        RECT 2547.315 14.090 2547.645 14.105 ;
        RECT 2621.145 14.090 2621.475 14.105 ;
        RECT 2547.315 13.790 2562.810 14.090 ;
        RECT 2547.315 13.775 2547.645 13.790 ;
        RECT 2562.510 13.410 2562.810 13.790 ;
        RECT 2586.430 13.790 2621.475 14.090 ;
        RECT 2586.430 13.410 2586.730 13.790 ;
        RECT 2621.145 13.775 2621.475 13.790 ;
        RECT 2562.510 13.110 2586.730 13.410 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.970 14.125 2564.110 15.300 ;
        RECT 2563.900 13.755 2564.180 14.125 ;
        RECT 2638.190 13.330 2638.470 13.445 ;
        RECT 2638.190 13.190 2639.320 13.330 ;
        RECT 2638.190 13.075 2638.470 13.190 ;
        RECT 2639.180 2.400 2639.320 13.190 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
      LAYER met3 ;
        RECT 2585.510 16.510 2638.250 16.810 ;
        RECT 2572.590 16.130 2572.970 16.140 ;
        RECT 2585.510 16.130 2585.810 16.510 ;
        RECT 2572.590 15.830 2585.810 16.130 ;
        RECT 2572.590 15.820 2572.970 15.830 ;
        RECT 2637.950 15.460 2638.250 16.510 ;
        RECT 2637.910 15.140 2638.290 15.460 ;
        RECT 2563.875 14.090 2564.205 14.105 ;
        RECT 2572.590 14.090 2572.970 14.100 ;
        RECT 2563.875 13.790 2572.970 14.090 ;
        RECT 2563.875 13.775 2564.205 13.790 ;
        RECT 2572.590 13.780 2572.970 13.790 ;
        RECT 2638.165 13.420 2638.495 13.425 ;
        RECT 2637.910 13.410 2638.495 13.420 ;
        RECT 2637.910 13.110 2638.720 13.410 ;
        RECT 2637.910 13.100 2638.495 13.110 ;
        RECT 2638.165 13.095 2638.495 13.100 ;
      LAYER met4 ;
        RECT 2572.615 15.815 2572.945 16.145 ;
        RECT 2572.630 14.105 2572.930 15.815 ;
        RECT 2637.935 15.135 2638.265 15.465 ;
        RECT 2572.615 13.775 2572.945 14.105 ;
        RECT 2637.950 13.425 2638.250 15.135 ;
        RECT 2637.935 13.095 2638.265 13.425 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2580.210 6.360 2580.530 6.420 ;
        RECT 2656.570 6.360 2656.890 6.420 ;
        RECT 2580.210 6.220 2656.890 6.360 ;
        RECT 2580.210 6.160 2580.530 6.220 ;
        RECT 2656.570 6.160 2656.890 6.220 ;
      LAYER met2 ;
        RECT 2580.530 14.010 2580.670 15.300 ;
        RECT 2580.300 13.870 2580.670 14.010 ;
        RECT 2580.300 6.450 2580.440 13.870 ;
        RECT 2580.240 6.130 2580.500 6.450 ;
        RECT 2656.600 6.130 2656.860 6.450 ;
        RECT 2656.660 2.400 2656.800 6.130 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.090 14.010 2597.230 15.300 ;
        RECT 2596.860 13.870 2597.230 14.010 ;
        RECT 2596.860 2.565 2597.000 13.870 ;
        RECT 2673.680 2.990 2674.740 3.130 ;
        RECT 2596.790 2.195 2597.070 2.565 ;
        RECT 2673.680 0.525 2673.820 2.990 ;
        RECT 2674.600 2.400 2674.740 2.990 ;
        RECT 2673.610 0.155 2673.890 0.525 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
      LAYER met3 ;
        RECT 2596.765 2.530 2597.095 2.545 ;
        RECT 2596.550 2.215 2597.095 2.530 ;
        RECT 2596.550 0.490 2596.850 2.215 ;
        RECT 2673.585 0.490 2673.915 0.505 ;
        RECT 2596.550 0.190 2673.915 0.490 ;
        RECT 2673.585 0.175 2673.915 0.190 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2613.790 0.920 2614.110 0.980 ;
        RECT 2691.070 0.920 2691.390 0.980 ;
        RECT 2613.790 0.780 2691.390 0.920 ;
        RECT 2613.790 0.720 2614.110 0.780 ;
        RECT 2691.070 0.720 2691.390 0.780 ;
      LAYER met2 ;
        RECT 2613.650 14.010 2613.790 15.300 ;
        RECT 2613.650 13.870 2614.020 14.010 ;
        RECT 2613.880 1.010 2614.020 13.870 ;
        RECT 2691.870 1.090 2692.430 2.400 ;
        RECT 2691.160 1.010 2692.430 1.090 ;
        RECT 2613.820 0.690 2614.080 1.010 ;
        RECT 2691.100 0.950 2692.430 1.010 ;
        RECT 2691.100 0.690 2691.360 0.950 ;
        RECT 2691.870 -4.800 2692.430 0.950 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.210 13.870 2630.350 15.300 ;
        RECT 2630.210 13.730 2630.580 13.870 ;
        RECT 2630.440 1.205 2630.580 13.730 ;
        RECT 2630.370 0.835 2630.650 1.205 ;
        RECT 2709.810 1.090 2710.370 2.400 ;
        RECT 2710.870 1.090 2711.150 1.205 ;
        RECT 2709.810 0.950 2711.150 1.090 ;
        RECT 2709.810 -4.800 2710.370 0.950 ;
        RECT 2710.870 0.835 2711.150 0.950 ;
      LAYER met3 ;
        RECT 2630.345 1.170 2630.675 1.185 ;
        RECT 2710.845 1.170 2711.175 1.185 ;
        RECT 2630.345 0.870 2711.175 1.170 ;
        RECT 2630.345 0.855 2630.675 0.870 ;
        RECT 2710.845 0.855 2711.175 0.870 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.770 14.805 2646.910 15.300 ;
        RECT 2646.700 14.435 2646.980 14.805 ;
        RECT 2726.510 12.650 2726.790 12.765 ;
        RECT 2726.510 12.510 2727.640 12.650 ;
        RECT 2726.510 12.395 2726.790 12.510 ;
        RECT 2727.500 2.400 2727.640 12.510 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
      LAYER met3 ;
        RECT 2726.230 18.170 2726.610 18.180 ;
        RECT 2653.590 17.870 2726.610 18.170 ;
        RECT 2646.675 14.770 2647.005 14.785 ;
        RECT 2653.590 14.770 2653.890 17.870 ;
        RECT 2726.230 17.860 2726.610 17.870 ;
        RECT 2646.675 14.470 2653.890 14.770 ;
        RECT 2646.675 14.455 2647.005 14.470 ;
        RECT 2726.485 12.740 2726.815 12.745 ;
        RECT 2726.230 12.730 2726.815 12.740 ;
        RECT 2726.230 12.430 2727.040 12.730 ;
        RECT 2726.230 12.420 2726.815 12.430 ;
        RECT 2726.485 12.415 2726.815 12.420 ;
      LAYER met4 ;
        RECT 2726.255 17.855 2726.585 18.185 ;
        RECT 2726.270 12.745 2726.570 17.855 ;
        RECT 2726.255 12.415 2726.585 12.745 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2663.470 1.600 2663.790 1.660 ;
        RECT 2743.510 1.600 2743.830 1.660 ;
        RECT 2663.470 1.460 2743.830 1.600 ;
        RECT 2663.470 1.400 2663.790 1.460 ;
        RECT 2743.510 1.400 2743.830 1.460 ;
      LAYER met2 ;
        RECT 2663.330 13.870 2663.470 15.300 ;
        RECT 2663.100 13.730 2663.470 13.870 ;
        RECT 2663.100 3.130 2663.240 13.730 ;
        RECT 2663.100 2.990 2663.700 3.130 ;
        RECT 2663.560 1.690 2663.700 2.990 ;
        RECT 2745.230 1.770 2745.790 2.400 ;
        RECT 2743.600 1.690 2745.790 1.770 ;
        RECT 2663.500 1.370 2663.760 1.690 ;
        RECT 2743.540 1.630 2745.790 1.690 ;
        RECT 2743.540 1.370 2743.800 1.630 ;
        RECT 2745.230 -4.800 2745.790 1.630 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.850 14.010 874.990 15.300 ;
        RECT 874.620 13.870 874.990 14.010 ;
        RECT 829.540 2.990 830.600 3.130 ;
        RECT 829.540 1.885 829.680 2.990 ;
        RECT 830.460 2.400 830.600 2.990 ;
        RECT 829.470 1.515 829.750 1.885 ;
        RECT 830.250 -4.800 830.810 2.400 ;
        RECT 874.620 1.885 874.760 13.870 ;
        RECT 874.550 1.515 874.830 1.885 ;
      LAYER met3 ;
        RECT 829.445 1.850 829.775 1.865 ;
        RECT 874.525 1.850 874.855 1.865 ;
        RECT 829.445 1.550 874.855 1.850 ;
        RECT 829.445 1.535 829.775 1.550 ;
        RECT 874.525 1.535 874.855 1.550 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2679.890 14.805 2680.030 15.300 ;
        RECT 2679.820 14.435 2680.100 14.805 ;
        RECT 2762.390 13.075 2762.670 13.445 ;
        RECT 2762.460 3.810 2762.600 13.075 ;
        RECT 2762.460 3.670 2763.520 3.810 ;
        RECT 2763.380 2.400 2763.520 3.670 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
      LAYER met3 ;
        RECT 2762.110 16.810 2762.490 16.820 ;
        RECT 2737.310 16.510 2762.490 16.810 ;
        RECT 2737.310 16.130 2737.610 16.510 ;
        RECT 2762.110 16.500 2762.490 16.510 ;
        RECT 2690.850 15.830 2737.610 16.130 ;
        RECT 2679.795 14.770 2680.125 14.785 ;
        RECT 2690.850 14.770 2691.150 15.830 ;
        RECT 2679.795 14.470 2691.150 14.770 ;
        RECT 2679.795 14.455 2680.125 14.470 ;
        RECT 2762.365 13.420 2762.695 13.425 ;
        RECT 2762.110 13.410 2762.695 13.420 ;
        RECT 2762.110 13.110 2762.920 13.410 ;
        RECT 2762.110 13.100 2762.695 13.110 ;
        RECT 2762.365 13.095 2762.695 13.100 ;
      LAYER met4 ;
        RECT 2762.135 16.495 2762.465 16.825 ;
        RECT 2762.150 13.425 2762.450 16.495 ;
        RECT 2762.135 13.095 2762.465 13.425 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2696.590 2.280 2696.910 2.340 ;
        RECT 2781.690 2.280 2782.010 2.340 ;
        RECT 2696.590 2.140 2782.010 2.280 ;
        RECT 2696.590 2.080 2696.910 2.140 ;
        RECT 2781.690 2.080 2782.010 2.140 ;
      LAYER met2 ;
        RECT 2696.450 14.010 2696.590 15.300 ;
        RECT 2696.450 13.870 2696.820 14.010 ;
        RECT 2696.680 2.370 2696.820 13.870 ;
        RECT 2696.620 2.050 2696.880 2.370 ;
        RECT 2780.650 1.770 2781.210 2.400 ;
        RECT 2781.720 2.050 2781.980 2.370 ;
        RECT 2781.780 1.770 2781.920 2.050 ;
        RECT 2780.650 1.630 2781.920 1.770 ;
        RECT 2780.650 -4.800 2781.210 1.630 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2713.010 14.125 2713.150 15.300 ;
        RECT 2712.940 13.755 2713.220 14.125 ;
        RECT 2796.430 12.650 2796.710 12.765 ;
        RECT 2796.430 12.510 2797.100 12.650 ;
        RECT 2796.430 12.395 2796.710 12.510 ;
        RECT 2796.960 1.770 2797.100 12.510 ;
        RECT 2798.590 1.770 2799.150 2.400 ;
        RECT 2796.960 1.630 2799.150 1.770 ;
        RECT 2798.590 -4.800 2799.150 1.630 ;
      LAYER met3 ;
        RECT 2712.915 14.090 2713.245 14.105 ;
        RECT 2712.915 13.790 2791.890 14.090 ;
        RECT 2712.915 13.775 2713.245 13.790 ;
        RECT 2791.590 12.730 2791.890 13.790 ;
        RECT 2796.405 12.730 2796.735 12.745 ;
        RECT 2791.590 12.430 2796.735 12.730 ;
        RECT 2796.405 12.415 2796.735 12.430 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2729.570 13.870 2729.710 15.300 ;
        RECT 2729.570 13.730 2729.940 13.870 ;
        RECT 2729.800 3.925 2729.940 13.730 ;
        RECT 2729.730 3.555 2730.010 3.925 ;
        RECT 2816.210 3.555 2816.490 3.925 ;
        RECT 2816.280 2.400 2816.420 3.555 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
      LAYER met3 ;
        RECT 2729.705 3.890 2730.035 3.905 ;
        RECT 2816.185 3.890 2816.515 3.905 ;
        RECT 2729.705 3.590 2816.515 3.890 ;
        RECT 2729.705 3.575 2730.035 3.590 ;
        RECT 2816.185 3.575 2816.515 3.590 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2745.810 5.680 2746.130 5.740 ;
        RECT 2834.130 5.680 2834.450 5.740 ;
        RECT 2745.810 5.540 2834.450 5.680 ;
        RECT 2745.810 5.480 2746.130 5.540 ;
        RECT 2834.130 5.480 2834.450 5.540 ;
      LAYER met2 ;
        RECT 2746.130 13.870 2746.270 15.300 ;
        RECT 2745.900 13.730 2746.270 13.870 ;
        RECT 2745.900 5.770 2746.040 13.730 ;
        RECT 2745.840 5.450 2746.100 5.770 ;
        RECT 2834.160 5.450 2834.420 5.770 ;
        RECT 2834.220 2.400 2834.360 5.450 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2762.690 13.870 2762.830 15.300 ;
        RECT 2762.690 13.730 2763.060 13.870 ;
        RECT 2762.920 4.605 2763.060 13.730 ;
        RECT 2762.850 4.235 2763.130 4.605 ;
        RECT 2851.630 4.235 2851.910 4.605 ;
        RECT 2851.700 2.400 2851.840 4.235 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
      LAYER met3 ;
        RECT 2762.825 4.570 2763.155 4.585 ;
        RECT 2851.605 4.570 2851.935 4.585 ;
        RECT 2762.825 4.270 2851.935 4.570 ;
        RECT 2762.825 4.255 2763.155 4.270 ;
        RECT 2851.605 4.255 2851.935 4.270 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2779.390 6.020 2779.710 6.080 ;
        RECT 2866.790 6.020 2867.110 6.080 ;
        RECT 2779.390 5.880 2867.110 6.020 ;
        RECT 2779.390 5.820 2779.710 5.880 ;
        RECT 2866.790 5.820 2867.110 5.880 ;
      LAYER met2 ;
        RECT 2779.250 14.010 2779.390 15.300 ;
        RECT 2779.250 13.870 2779.620 14.010 ;
        RECT 2779.480 6.110 2779.620 13.870 ;
        RECT 2779.420 5.790 2779.680 6.110 ;
        RECT 2866.820 5.790 2867.080 6.110 ;
        RECT 2866.880 1.770 2867.020 5.790 ;
        RECT 2869.430 1.770 2869.990 2.400 ;
        RECT 2866.880 1.630 2869.990 1.770 ;
        RECT 2869.430 -4.800 2869.990 1.630 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2795.810 14.010 2795.950 15.300 ;
        RECT 2795.810 13.870 2796.180 14.010 ;
        RECT 2796.040 2.565 2796.180 13.870 ;
        RECT 2795.970 2.195 2796.250 2.565 ;
        RECT 2885.670 2.195 2885.950 2.565 ;
        RECT 2885.740 1.770 2885.880 2.195 ;
        RECT 2886.910 1.770 2887.470 2.400 ;
        RECT 2885.740 1.630 2887.470 1.770 ;
        RECT 2886.910 -4.800 2887.470 1.630 ;
      LAYER met3 ;
        RECT 2795.945 2.530 2796.275 2.545 ;
        RECT 2885.645 2.530 2885.975 2.545 ;
        RECT 2795.945 2.230 2885.975 2.530 ;
        RECT 2795.945 2.215 2796.275 2.230 ;
        RECT 2885.645 2.215 2885.975 2.230 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 847.850 14.520 848.170 14.580 ;
        RECT 891.320 14.520 891.640 14.580 ;
        RECT 847.850 14.380 891.640 14.520 ;
        RECT 847.850 14.320 848.170 14.380 ;
        RECT 891.320 14.320 891.640 14.380 ;
      LAYER met2 ;
        RECT 891.410 14.610 891.550 15.300 ;
        RECT 847.880 14.290 848.140 14.610 ;
        RECT 891.350 14.290 891.610 14.610 ;
        RECT 847.940 2.400 848.080 14.290 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.970 14.010 908.110 15.300 ;
        RECT 907.740 13.870 908.110 14.010 ;
        RECT 907.740 3.245 907.880 13.870 ;
        RECT 865.810 2.875 866.090 3.245 ;
        RECT 907.670 2.875 907.950 3.245 ;
        RECT 865.880 2.400 866.020 2.875 ;
        RECT 865.670 -4.800 866.230 2.400 ;
      LAYER met3 ;
        RECT 865.785 3.210 866.115 3.225 ;
        RECT 907.645 3.210 907.975 3.225 ;
        RECT 865.785 2.910 907.975 3.210 ;
        RECT 865.785 2.895 866.115 2.910 ;
        RECT 907.645 2.895 907.975 2.910 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.530 14.010 924.670 15.300 ;
        RECT 924.300 13.870 924.670 14.010 ;
        RECT 924.300 3.245 924.440 13.870 ;
        RECT 883.360 2.990 884.420 3.130 ;
        RECT 883.360 2.400 883.500 2.990 ;
        RECT 883.150 -4.800 883.710 2.400 ;
        RECT 884.280 1.885 884.420 2.990 ;
        RECT 924.230 2.875 924.510 3.245 ;
        RECT 884.210 1.515 884.490 1.885 ;
      LAYER met3 ;
        RECT 924.205 3.210 924.535 3.225 ;
        RECT 913.870 2.910 924.535 3.210 ;
        RECT 884.185 1.850 884.515 1.865 ;
        RECT 913.870 1.850 914.170 2.910 ;
        RECT 924.205 2.895 924.535 2.910 ;
        RECT 884.185 1.550 914.170 1.850 ;
        RECT 884.185 1.535 884.515 1.550 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.090 14.010 941.230 15.300 ;
        RECT 940.860 13.870 941.230 14.010 ;
        RECT 940.860 10.045 941.000 13.870 ;
        RECT 901.230 9.675 901.510 10.045 ;
        RECT 940.790 9.675 941.070 10.045 ;
        RECT 901.300 2.400 901.440 9.675 ;
        RECT 901.090 -4.800 901.650 2.400 ;
      LAYER met3 ;
        RECT 901.205 10.010 901.535 10.025 ;
        RECT 940.765 10.010 941.095 10.025 ;
        RECT 901.205 9.710 941.095 10.010 ;
        RECT 901.205 9.695 901.535 9.710 ;
        RECT 940.765 9.695 941.095 9.710 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.650 14.010 957.790 15.300 ;
        RECT 957.420 13.870 957.790 14.010 ;
        RECT 957.420 5.965 957.560 13.870 ;
        RECT 918.710 5.595 918.990 5.965 ;
        RECT 957.350 5.595 957.630 5.965 ;
        RECT 918.780 2.400 918.920 5.595 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER met3 ;
        RECT 918.685 5.930 919.015 5.945 ;
        RECT 957.325 5.930 957.655 5.945 ;
        RECT 918.685 5.630 957.655 5.930 ;
        RECT 918.685 5.615 919.015 5.630 ;
        RECT 957.325 5.615 957.655 5.630 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.210 14.010 974.350 15.300 ;
        RECT 973.980 13.870 974.350 14.010 ;
        RECT 935.730 0.410 936.010 0.525 ;
        RECT 936.510 0.410 937.070 2.400 ;
        RECT 973.980 0.525 974.120 13.870 ;
        RECT 935.730 0.270 937.070 0.410 ;
        RECT 935.730 0.155 936.010 0.270 ;
        RECT 936.510 -4.800 937.070 0.270 ;
        RECT 973.910 0.155 974.190 0.525 ;
      LAYER met3 ;
        RECT 935.705 0.490 936.035 0.505 ;
        RECT 973.885 0.490 974.215 0.505 ;
        RECT 935.705 0.190 974.215 0.490 ;
        RECT 935.705 0.175 936.035 0.190 ;
        RECT 973.885 0.175 974.215 0.190 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.770 14.010 990.910 15.300 ;
        RECT 990.540 13.870 990.910 14.010 ;
        RECT 990.540 3.925 990.680 13.870 ;
        RECT 954.130 3.555 954.410 3.925 ;
        RECT 990.470 3.555 990.750 3.925 ;
        RECT 954.200 2.400 954.340 3.555 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER met3 ;
        RECT 954.105 3.890 954.435 3.905 ;
        RECT 990.445 3.890 990.775 3.905 ;
        RECT 954.105 3.590 990.775 3.890 ;
        RECT 954.105 3.575 954.435 3.590 ;
        RECT 990.445 3.575 990.775 3.590 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.330 14.010 1007.470 15.300 ;
        RECT 1007.100 13.870 1007.470 14.010 ;
        RECT 1007.100 5.965 1007.240 13.870 ;
        RECT 972.070 5.595 972.350 5.965 ;
        RECT 1007.030 5.595 1007.310 5.965 ;
        RECT 972.140 2.400 972.280 5.595 ;
        RECT 971.930 -4.800 972.490 2.400 ;
      LAYER met3 ;
        RECT 972.045 5.930 972.375 5.945 ;
        RECT 1007.005 5.930 1007.335 5.945 ;
        RECT 972.045 5.630 1007.335 5.930 ;
        RECT 972.045 5.615 972.375 5.630 ;
        RECT 1007.005 5.615 1007.335 5.630 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.250 14.010 709.390 15.300 ;
        RECT 709.020 13.870 709.390 14.010 ;
        RECT 709.020 5.285 709.160 13.870 ;
        RECT 663.870 4.915 664.150 5.285 ;
        RECT 708.950 4.915 709.230 5.285 ;
        RECT 663.940 3.245 664.080 4.915 ;
        RECT 652.830 2.875 653.110 3.245 ;
        RECT 663.870 2.875 664.150 3.245 ;
        RECT 652.900 2.400 653.040 2.875 ;
        RECT 652.690 -4.800 653.250 2.400 ;
      LAYER met3 ;
        RECT 663.845 5.250 664.175 5.265 ;
        RECT 708.925 5.250 709.255 5.265 ;
        RECT 663.845 4.950 709.255 5.250 ;
        RECT 663.845 4.935 664.175 4.950 ;
        RECT 708.925 4.935 709.255 4.950 ;
        RECT 652.805 3.210 653.135 3.225 ;
        RECT 663.845 3.210 664.175 3.225 ;
        RECT 652.805 2.910 664.175 3.210 ;
        RECT 652.805 2.895 653.135 2.910 ;
        RECT 663.845 2.895 664.175 2.910 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.890 14.010 1024.030 15.300 ;
        RECT 1023.660 13.870 1024.030 14.010 ;
        RECT 989.410 1.770 989.970 2.400 ;
        RECT 1023.660 1.885 1023.800 13.870 ;
        RECT 991.850 1.770 992.130 1.885 ;
        RECT 989.410 1.630 992.130 1.770 ;
        RECT 989.410 -4.800 989.970 1.630 ;
        RECT 991.850 1.515 992.130 1.630 ;
        RECT 1023.590 1.515 1023.870 1.885 ;
      LAYER met3 ;
        RECT 991.825 1.850 992.155 1.865 ;
        RECT 1023.565 1.850 1023.895 1.865 ;
        RECT 991.825 1.550 1023.895 1.850 ;
        RECT 991.825 1.535 992.155 1.550 ;
        RECT 1023.565 1.535 1023.895 1.550 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.450 14.010 1040.590 15.300 ;
        RECT 1040.220 13.870 1040.590 14.010 ;
        RECT 1040.220 7.325 1040.360 13.870 ;
        RECT 1007.490 6.955 1007.770 7.325 ;
        RECT 1040.150 6.955 1040.430 7.325 ;
        RECT 1007.560 2.400 1007.700 6.955 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER met3 ;
        RECT 1007.465 7.290 1007.795 7.305 ;
        RECT 1040.125 7.290 1040.455 7.305 ;
        RECT 1007.465 6.990 1040.455 7.290 ;
        RECT 1007.465 6.975 1007.795 6.990 ;
        RECT 1040.125 6.975 1040.455 6.990 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.010 14.010 1057.150 15.300 ;
        RECT 1056.780 13.870 1057.150 14.010 ;
        RECT 1056.780 6.645 1056.920 13.870 ;
        RECT 1025.430 6.275 1025.710 6.645 ;
        RECT 1056.710 6.275 1056.990 6.645 ;
        RECT 1025.500 2.400 1025.640 6.275 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
      LAYER met3 ;
        RECT 1025.405 6.610 1025.735 6.625 ;
        RECT 1056.685 6.610 1057.015 6.625 ;
        RECT 1025.405 6.310 1057.015 6.610 ;
        RECT 1025.405 6.295 1025.735 6.310 ;
        RECT 1056.685 6.295 1057.015 6.310 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.570 14.010 1073.710 15.300 ;
        RECT 1073.340 13.870 1073.710 14.010 ;
        RECT 1073.340 10.045 1073.480 13.870 ;
        RECT 1042.910 9.675 1043.190 10.045 ;
        RECT 1073.270 9.675 1073.550 10.045 ;
        RECT 1042.980 2.400 1043.120 9.675 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
      LAYER met3 ;
        RECT 1042.885 10.010 1043.215 10.025 ;
        RECT 1073.245 10.010 1073.575 10.025 ;
        RECT 1042.885 9.710 1073.575 10.010 ;
        RECT 1042.885 9.695 1043.215 9.710 ;
        RECT 1073.245 9.695 1073.575 9.710 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.130 14.010 1090.270 15.300 ;
        RECT 1089.900 13.870 1090.270 14.010 ;
        RECT 1089.900 9.365 1090.040 13.870 ;
        RECT 1060.850 8.995 1061.130 9.365 ;
        RECT 1089.830 8.995 1090.110 9.365 ;
        RECT 1060.920 2.400 1061.060 8.995 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
      LAYER met3 ;
        RECT 1060.825 9.330 1061.155 9.345 ;
        RECT 1089.805 9.330 1090.135 9.345 ;
        RECT 1060.825 9.030 1090.135 9.330 ;
        RECT 1060.825 9.015 1061.155 9.030 ;
        RECT 1089.805 9.015 1090.135 9.030 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.690 14.010 1106.830 15.300 ;
        RECT 1106.460 13.870 1106.830 14.010 ;
        RECT 1106.460 8.005 1106.600 13.870 ;
        RECT 1078.330 7.635 1078.610 8.005 ;
        RECT 1106.390 7.635 1106.670 8.005 ;
        RECT 1078.400 2.400 1078.540 7.635 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
      LAYER met3 ;
        RECT 1078.305 7.970 1078.635 7.985 ;
        RECT 1106.365 7.970 1106.695 7.985 ;
        RECT 1078.305 7.670 1106.695 7.970 ;
        RECT 1078.305 7.655 1078.635 7.670 ;
        RECT 1106.365 7.655 1106.695 7.670 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.250 14.010 1123.390 15.300 ;
        RECT 1123.020 13.870 1123.390 14.010 ;
        RECT 1123.020 11.405 1123.160 13.870 ;
        RECT 1096.270 11.035 1096.550 11.405 ;
        RECT 1122.950 11.035 1123.230 11.405 ;
        RECT 1096.340 2.400 1096.480 11.035 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
      LAYER met3 ;
        RECT 1096.245 11.370 1096.575 11.385 ;
        RECT 1122.925 11.370 1123.255 11.385 ;
        RECT 1096.245 11.070 1123.255 11.370 ;
        RECT 1096.245 11.055 1096.575 11.070 ;
        RECT 1122.925 11.055 1123.255 11.070 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.810 14.010 1139.950 15.300 ;
        RECT 1139.580 13.870 1139.950 14.010 ;
        RECT 1139.580 8.685 1139.720 13.870 ;
        RECT 1113.750 8.315 1114.030 8.685 ;
        RECT 1139.510 8.315 1139.790 8.685 ;
        RECT 1113.820 2.400 1113.960 8.315 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
      LAYER met3 ;
        RECT 1113.725 8.650 1114.055 8.665 ;
        RECT 1139.485 8.650 1139.815 8.665 ;
        RECT 1113.725 8.350 1139.815 8.650 ;
        RECT 1113.725 8.335 1114.055 8.350 ;
        RECT 1139.485 8.335 1139.815 8.350 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.370 14.010 1156.510 15.300 ;
        RECT 1156.140 13.870 1156.510 14.010 ;
        RECT 1156.140 8.005 1156.280 13.870 ;
        RECT 1131.690 7.635 1131.970 8.005 ;
        RECT 1156.070 7.635 1156.350 8.005 ;
        RECT 1131.760 2.400 1131.900 7.635 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
      LAYER met3 ;
        RECT 1131.665 7.970 1131.995 7.985 ;
        RECT 1156.045 7.970 1156.375 7.985 ;
        RECT 1131.665 7.670 1156.375 7.970 ;
        RECT 1131.665 7.655 1131.995 7.670 ;
        RECT 1156.045 7.655 1156.375 7.670 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.930 14.010 1173.070 15.300 ;
        RECT 1172.700 13.870 1173.070 14.010 ;
        RECT 1172.700 10.725 1172.840 13.870 ;
        RECT 1149.170 10.355 1149.450 10.725 ;
        RECT 1172.630 10.355 1172.910 10.725 ;
        RECT 1149.240 2.400 1149.380 10.355 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
      LAYER met3 ;
        RECT 1149.145 10.690 1149.475 10.705 ;
        RECT 1172.605 10.690 1172.935 10.705 ;
        RECT 1149.145 10.390 1172.935 10.690 ;
        RECT 1149.145 10.375 1149.475 10.390 ;
        RECT 1172.605 10.375 1172.935 10.390 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 671.670 14.520 671.990 14.580 ;
        RECT 725.720 14.520 726.040 14.580 ;
        RECT 671.670 14.380 726.040 14.520 ;
        RECT 671.670 14.320 671.990 14.380 ;
        RECT 725.720 14.320 726.040 14.380 ;
      LAYER met2 ;
        RECT 725.810 14.610 725.950 15.300 ;
        RECT 671.700 14.290 671.960 14.610 ;
        RECT 725.750 14.290 726.010 14.610 ;
        RECT 671.760 7.210 671.900 14.290 ;
        RECT 670.840 7.070 671.900 7.210 ;
        RECT 670.840 2.400 670.980 7.070 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.490 14.010 1189.630 15.300 ;
        RECT 1189.260 13.870 1189.630 14.010 ;
        RECT 1189.260 9.365 1189.400 13.870 ;
        RECT 1167.110 8.995 1167.390 9.365 ;
        RECT 1189.190 8.995 1189.470 9.365 ;
        RECT 1167.180 2.400 1167.320 8.995 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
      LAYER met3 ;
        RECT 1167.085 9.330 1167.415 9.345 ;
        RECT 1189.165 9.330 1189.495 9.345 ;
        RECT 1167.085 9.030 1189.495 9.330 ;
        RECT 1167.085 9.015 1167.415 9.030 ;
        RECT 1189.165 9.015 1189.495 9.030 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.050 14.010 1206.190 15.300 ;
        RECT 1205.820 13.870 1206.190 14.010 ;
        RECT 1205.820 8.005 1205.960 13.870 ;
        RECT 1185.050 7.635 1185.330 8.005 ;
        RECT 1205.750 7.635 1206.030 8.005 ;
        RECT 1185.120 2.400 1185.260 7.635 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
      LAYER met3 ;
        RECT 1185.025 7.970 1185.355 7.985 ;
        RECT 1205.725 7.970 1206.055 7.985 ;
        RECT 1185.025 7.670 1206.055 7.970 ;
        RECT 1185.025 7.655 1185.355 7.670 ;
        RECT 1205.725 7.655 1206.055 7.670 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.610 14.010 1222.750 15.300 ;
        RECT 1222.380 13.870 1222.750 14.010 ;
        RECT 1222.380 7.325 1222.520 13.870 ;
        RECT 1202.530 6.955 1202.810 7.325 ;
        RECT 1222.310 6.955 1222.590 7.325 ;
        RECT 1202.600 2.400 1202.740 6.955 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
      LAYER met3 ;
        RECT 1202.505 7.290 1202.835 7.305 ;
        RECT 1222.285 7.290 1222.615 7.305 ;
        RECT 1202.505 6.990 1222.615 7.290 ;
        RECT 1202.505 6.975 1202.835 6.990 ;
        RECT 1222.285 6.975 1222.615 6.990 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.170 14.010 1239.310 15.300 ;
        RECT 1238.940 13.870 1239.310 14.010 ;
        RECT 1238.940 8.005 1239.080 13.870 ;
        RECT 1220.470 7.635 1220.750 8.005 ;
        RECT 1238.870 7.635 1239.150 8.005 ;
        RECT 1220.540 2.400 1220.680 7.635 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
      LAYER met3 ;
        RECT 1220.445 7.970 1220.775 7.985 ;
        RECT 1238.845 7.970 1239.175 7.985 ;
        RECT 1220.445 7.670 1239.175 7.970 ;
        RECT 1220.445 7.655 1220.775 7.670 ;
        RECT 1238.845 7.655 1239.175 7.670 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.730 14.010 1255.870 15.300 ;
        RECT 1255.500 13.870 1255.870 14.010 ;
        RECT 1255.500 9.365 1255.640 13.870 ;
        RECT 1237.950 8.995 1238.230 9.365 ;
        RECT 1255.430 8.995 1255.710 9.365 ;
        RECT 1238.020 2.400 1238.160 8.995 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
      LAYER met3 ;
        RECT 1237.925 9.330 1238.255 9.345 ;
        RECT 1255.405 9.330 1255.735 9.345 ;
        RECT 1237.925 9.030 1255.735 9.330 ;
        RECT 1237.925 9.015 1238.255 9.030 ;
        RECT 1255.405 9.015 1255.735 9.030 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.290 14.010 1272.430 15.300 ;
        RECT 1272.060 13.870 1272.430 14.010 ;
        RECT 1272.060 8.685 1272.200 13.870 ;
        RECT 1255.890 8.315 1256.170 8.685 ;
        RECT 1271.990 8.315 1272.270 8.685 ;
        RECT 1255.960 2.400 1256.100 8.315 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
      LAYER met3 ;
        RECT 1255.865 8.650 1256.195 8.665 ;
        RECT 1271.965 8.650 1272.295 8.665 ;
        RECT 1255.865 8.350 1272.295 8.650 ;
        RECT 1255.865 8.335 1256.195 8.350 ;
        RECT 1271.965 8.335 1272.295 8.350 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.850 14.010 1288.990 15.300 ;
        RECT 1288.620 13.870 1288.990 14.010 ;
        RECT 1288.620 8.685 1288.760 13.870 ;
        RECT 1273.370 8.315 1273.650 8.685 ;
        RECT 1288.550 8.315 1288.830 8.685 ;
        RECT 1273.440 2.400 1273.580 8.315 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
      LAYER met3 ;
        RECT 1273.345 8.650 1273.675 8.665 ;
        RECT 1288.525 8.650 1288.855 8.665 ;
        RECT 1273.345 8.350 1288.855 8.650 ;
        RECT 1273.345 8.335 1273.675 8.350 ;
        RECT 1288.525 8.335 1288.855 8.350 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.410 14.010 1305.550 15.300 ;
        RECT 1305.180 13.870 1305.550 14.010 ;
        RECT 1305.180 8.685 1305.320 13.870 ;
        RECT 1291.310 8.315 1291.590 8.685 ;
        RECT 1305.110 8.315 1305.390 8.685 ;
        RECT 1291.380 2.400 1291.520 8.315 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
      LAYER met3 ;
        RECT 1291.285 8.650 1291.615 8.665 ;
        RECT 1305.085 8.650 1305.415 8.665 ;
        RECT 1291.285 8.350 1305.415 8.650 ;
        RECT 1291.285 8.335 1291.615 8.350 ;
        RECT 1305.085 8.335 1305.415 8.350 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.970 14.010 1322.110 15.300 ;
        RECT 1321.740 13.870 1322.110 14.010 ;
        RECT 1321.740 8.685 1321.880 13.870 ;
        RECT 1308.790 8.315 1309.070 8.685 ;
        RECT 1321.670 8.315 1321.950 8.685 ;
        RECT 1308.860 2.400 1309.000 8.315 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
      LAYER met3 ;
        RECT 1308.765 8.650 1309.095 8.665 ;
        RECT 1321.645 8.650 1321.975 8.665 ;
        RECT 1308.765 8.350 1321.975 8.650 ;
        RECT 1308.765 8.335 1309.095 8.350 ;
        RECT 1321.645 8.335 1321.975 8.350 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.530 14.010 1338.670 15.300 ;
        RECT 1338.300 13.870 1338.670 14.010 ;
        RECT 1338.300 5.285 1338.440 13.870 ;
        RECT 1326.730 4.915 1327.010 5.285 ;
        RECT 1338.230 4.915 1338.510 5.285 ;
        RECT 1326.800 2.400 1326.940 4.915 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
      LAYER met3 ;
        RECT 1326.705 5.250 1327.035 5.265 ;
        RECT 1338.205 5.250 1338.535 5.265 ;
        RECT 1326.705 4.950 1338.535 5.250 ;
        RECT 1326.705 4.935 1327.035 4.950 ;
        RECT 1338.205 4.935 1338.535 4.950 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.370 14.010 742.510 15.300 ;
        RECT 742.370 13.870 742.740 14.010 ;
        RECT 742.600 2.565 742.740 13.870 ;
        RECT 687.330 1.090 687.610 1.205 ;
        RECT 688.110 1.090 688.670 2.400 ;
        RECT 742.530 2.195 742.810 2.565 ;
        RECT 687.330 0.950 688.670 1.090 ;
        RECT 687.330 0.835 687.610 0.950 ;
        RECT 688.110 -4.800 688.670 0.950 ;
      LAYER met3 ;
        RECT 742.505 2.530 742.835 2.545 ;
        RECT 742.505 2.215 743.050 2.530 ;
        RECT 687.305 1.170 687.635 1.185 ;
        RECT 742.750 1.170 743.050 2.215 ;
        RECT 687.305 0.870 743.050 1.170 ;
        RECT 687.305 0.855 687.635 0.870 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.090 14.010 1355.230 15.300 ;
        RECT 1354.860 13.870 1355.230 14.010 ;
        RECT 1354.860 7.325 1355.000 13.870 ;
        RECT 1344.210 6.955 1344.490 7.325 ;
        RECT 1354.790 6.955 1355.070 7.325 ;
        RECT 1344.280 2.400 1344.420 6.955 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
      LAYER met3 ;
        RECT 1344.185 7.290 1344.515 7.305 ;
        RECT 1354.765 7.290 1355.095 7.305 ;
        RECT 1344.185 6.990 1355.095 7.290 ;
        RECT 1344.185 6.975 1344.515 6.990 ;
        RECT 1354.765 6.975 1355.095 6.990 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.650 14.010 1371.790 15.300 ;
        RECT 1371.420 13.870 1371.790 14.010 ;
        RECT 1371.420 5.965 1371.560 13.870 ;
        RECT 1362.150 5.595 1362.430 5.965 ;
        RECT 1371.350 5.595 1371.630 5.965 ;
        RECT 1362.220 2.400 1362.360 5.595 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
      LAYER met3 ;
        RECT 1362.125 5.930 1362.455 5.945 ;
        RECT 1371.325 5.930 1371.655 5.945 ;
        RECT 1362.125 5.630 1371.655 5.930 ;
        RECT 1362.125 5.615 1362.455 5.630 ;
        RECT 1371.325 5.615 1371.655 5.630 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.210 14.010 1388.350 15.300 ;
        RECT 1387.980 13.870 1388.350 14.010 ;
        RECT 1387.980 6.645 1388.120 13.870 ;
        RECT 1380.090 6.275 1380.370 6.645 ;
        RECT 1387.910 6.275 1388.190 6.645 ;
        RECT 1380.160 2.400 1380.300 6.275 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
      LAYER met3 ;
        RECT 1380.065 6.610 1380.395 6.625 ;
        RECT 1387.885 6.610 1388.215 6.625 ;
        RECT 1380.065 6.310 1388.215 6.610 ;
        RECT 1380.065 6.295 1380.395 6.310 ;
        RECT 1387.885 6.295 1388.215 6.310 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.770 14.010 1404.910 15.300 ;
        RECT 1404.540 13.870 1404.910 14.010 ;
        RECT 1404.540 6.645 1404.680 13.870 ;
        RECT 1397.570 6.275 1397.850 6.645 ;
        RECT 1404.470 6.275 1404.750 6.645 ;
        RECT 1397.640 2.400 1397.780 6.275 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
      LAYER met3 ;
        RECT 1397.545 6.610 1397.875 6.625 ;
        RECT 1404.445 6.610 1404.775 6.625 ;
        RECT 1397.545 6.310 1404.775 6.610 ;
        RECT 1397.545 6.295 1397.875 6.310 ;
        RECT 1404.445 6.295 1404.775 6.310 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.330 14.690 1421.470 15.300 ;
        RECT 1416.500 14.550 1421.470 14.690 ;
        RECT 1416.500 5.850 1416.640 14.550 ;
        RECT 1415.580 5.710 1416.640 5.850 ;
        RECT 1415.580 2.400 1415.720 5.710 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.890 14.010 1438.030 15.300 ;
        RECT 1437.660 13.870 1438.030 14.010 ;
        RECT 1437.660 6.645 1437.800 13.870 ;
        RECT 1432.990 6.275 1433.270 6.645 ;
        RECT 1437.590 6.275 1437.870 6.645 ;
        RECT 1433.060 2.400 1433.200 6.275 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
      LAYER met3 ;
        RECT 1432.965 6.610 1433.295 6.625 ;
        RECT 1437.565 6.610 1437.895 6.625 ;
        RECT 1432.965 6.310 1437.895 6.610 ;
        RECT 1432.965 6.295 1433.295 6.310 ;
        RECT 1437.565 6.295 1437.895 6.310 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.450 14.010 1454.590 15.300 ;
        RECT 1451.000 13.870 1454.590 14.010 ;
        RECT 1451.000 2.400 1451.140 13.870 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.010 14.010 1471.150 15.300 ;
        RECT 1468.480 13.870 1471.150 14.010 ;
        RECT 1468.480 2.400 1468.620 13.870 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.570 14.010 1487.710 15.300 ;
        RECT 1487.340 13.870 1487.710 14.010 ;
        RECT 1486.210 1.770 1486.770 2.400 ;
        RECT 1487.340 1.770 1487.480 13.870 ;
        RECT 1486.210 1.630 1487.480 1.770 ;
        RECT 1486.210 -4.800 1486.770 1.630 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.130 14.010 1504.270 15.300 ;
        RECT 1503.900 13.870 1504.270 14.010 ;
        RECT 1503.900 2.400 1504.040 13.870 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.930 14.010 759.070 15.300 ;
        RECT 758.700 13.870 759.070 14.010 ;
        RECT 758.700 11.405 758.840 13.870 ;
        RECT 706.190 11.035 706.470 11.405 ;
        RECT 758.630 11.035 758.910 11.405 ;
        RECT 706.260 2.400 706.400 11.035 ;
        RECT 706.050 -4.800 706.610 2.400 ;
      LAYER met3 ;
        RECT 706.165 11.370 706.495 11.385 ;
        RECT 758.605 11.370 758.935 11.385 ;
        RECT 706.165 11.070 758.935 11.370 ;
        RECT 706.165 11.055 706.495 11.070 ;
        RECT 758.605 11.055 758.935 11.070 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.690 14.010 1520.830 15.300 ;
        RECT 1520.690 13.870 1521.060 14.010 ;
        RECT 1520.920 1.770 1521.060 13.870 ;
        RECT 1521.630 1.770 1522.190 2.400 ;
        RECT 1520.920 1.630 1522.190 1.770 ;
        RECT 1521.630 -4.800 1522.190 1.630 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.250 14.010 1537.390 15.300 ;
        RECT 1537.250 13.870 1539.920 14.010 ;
        RECT 1539.780 2.400 1539.920 13.870 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.810 14.010 1553.950 15.300 ;
        RECT 1553.810 13.870 1557.400 14.010 ;
        RECT 1557.260 2.400 1557.400 13.870 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.370 14.010 1570.510 15.300 ;
        RECT 1570.370 13.870 1570.740 14.010 ;
        RECT 1570.600 6.645 1570.740 13.870 ;
        RECT 1570.530 6.275 1570.810 6.645 ;
        RECT 1575.130 6.275 1575.410 6.645 ;
        RECT 1575.200 2.400 1575.340 6.275 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
      LAYER met3 ;
        RECT 1570.505 6.610 1570.835 6.625 ;
        RECT 1575.105 6.610 1575.435 6.625 ;
        RECT 1570.505 6.310 1575.435 6.610 ;
        RECT 1570.505 6.295 1570.835 6.310 ;
        RECT 1575.105 6.295 1575.435 6.310 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.930 14.690 1587.070 15.300 ;
        RECT 1586.930 14.550 1587.300 14.690 ;
        RECT 1587.160 6.645 1587.300 14.550 ;
        RECT 1587.090 6.275 1587.370 6.645 ;
        RECT 1592.610 6.275 1592.890 6.645 ;
        RECT 1592.680 2.400 1592.820 6.275 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
      LAYER met3 ;
        RECT 1587.065 6.610 1587.395 6.625 ;
        RECT 1592.585 6.610 1592.915 6.625 ;
        RECT 1587.065 6.310 1592.915 6.610 ;
        RECT 1587.065 6.295 1587.395 6.310 ;
        RECT 1592.585 6.295 1592.915 6.310 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.490 14.010 1603.630 15.300 ;
        RECT 1603.490 13.870 1603.860 14.010 ;
        RECT 1603.720 5.965 1603.860 13.870 ;
        RECT 1603.650 5.595 1603.930 5.965 ;
        RECT 1610.550 5.595 1610.830 5.965 ;
        RECT 1610.620 2.400 1610.760 5.595 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
      LAYER met3 ;
        RECT 1603.625 5.930 1603.955 5.945 ;
        RECT 1610.525 5.930 1610.855 5.945 ;
        RECT 1603.625 5.630 1610.855 5.930 ;
        RECT 1603.625 5.615 1603.955 5.630 ;
        RECT 1610.525 5.615 1610.855 5.630 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.050 14.010 1620.190 15.300 ;
        RECT 1620.050 13.870 1620.420 14.010 ;
        RECT 1620.280 5.965 1620.420 13.870 ;
        RECT 1620.210 5.595 1620.490 5.965 ;
        RECT 1628.030 5.595 1628.310 5.965 ;
        RECT 1628.100 2.400 1628.240 5.595 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
      LAYER met3 ;
        RECT 1620.185 5.930 1620.515 5.945 ;
        RECT 1628.005 5.930 1628.335 5.945 ;
        RECT 1620.185 5.630 1628.335 5.930 ;
        RECT 1620.185 5.615 1620.515 5.630 ;
        RECT 1628.005 5.615 1628.335 5.630 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.610 14.010 1636.750 15.300 ;
        RECT 1636.610 13.870 1636.980 14.010 ;
        RECT 1636.840 6.645 1636.980 13.870 ;
        RECT 1636.770 6.275 1637.050 6.645 ;
        RECT 1645.970 6.275 1646.250 6.645 ;
        RECT 1646.040 2.400 1646.180 6.275 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
      LAYER met3 ;
        RECT 1636.745 6.610 1637.075 6.625 ;
        RECT 1645.945 6.610 1646.275 6.625 ;
        RECT 1636.745 6.310 1646.275 6.610 ;
        RECT 1636.745 6.295 1637.075 6.310 ;
        RECT 1645.945 6.295 1646.275 6.310 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.170 14.010 1653.310 15.300 ;
        RECT 1653.170 13.870 1653.540 14.010 ;
        RECT 1653.400 5.965 1653.540 13.870 ;
        RECT 1653.330 5.595 1653.610 5.965 ;
        RECT 1663.450 5.595 1663.730 5.965 ;
        RECT 1663.520 2.400 1663.660 5.595 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
      LAYER met3 ;
        RECT 1653.305 5.930 1653.635 5.945 ;
        RECT 1663.425 5.930 1663.755 5.945 ;
        RECT 1653.305 5.630 1663.755 5.930 ;
        RECT 1653.305 5.615 1653.635 5.630 ;
        RECT 1663.425 5.615 1663.755 5.630 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.730 14.010 1669.870 15.300 ;
        RECT 1669.500 13.870 1669.870 14.010 ;
        RECT 1669.500 5.285 1669.640 13.870 ;
        RECT 1669.430 4.915 1669.710 5.285 ;
        RECT 1681.390 4.915 1681.670 5.285 ;
        RECT 1681.460 2.400 1681.600 4.915 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
      LAYER met3 ;
        RECT 1669.405 5.250 1669.735 5.265 ;
        RECT 1681.365 5.250 1681.695 5.265 ;
        RECT 1669.405 4.950 1681.695 5.250 ;
        RECT 1669.405 4.935 1669.735 4.950 ;
        RECT 1681.365 4.935 1681.695 4.950 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.570 0.920 724.890 0.980 ;
        RECT 775.170 0.920 775.490 0.980 ;
        RECT 724.570 0.780 775.490 0.920 ;
        RECT 724.570 0.720 724.890 0.780 ;
        RECT 775.170 0.720 775.490 0.780 ;
      LAYER met2 ;
        RECT 775.490 14.010 775.630 15.300 ;
        RECT 775.260 13.870 775.630 14.010 ;
        RECT 723.530 1.090 724.090 2.400 ;
        RECT 723.530 1.010 724.800 1.090 ;
        RECT 775.260 1.010 775.400 13.870 ;
        RECT 723.530 0.950 724.860 1.010 ;
        RECT 723.530 -4.800 724.090 0.950 ;
        RECT 724.600 0.690 724.860 0.950 ;
        RECT 775.200 0.690 775.460 1.010 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.290 14.010 1686.430 15.300 ;
        RECT 1686.290 13.870 1686.660 14.010 ;
        RECT 1686.520 5.285 1686.660 13.870 ;
        RECT 1686.450 4.915 1686.730 5.285 ;
        RECT 1699.330 4.915 1699.610 5.285 ;
        RECT 1699.400 2.400 1699.540 4.915 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
      LAYER met3 ;
        RECT 1686.425 5.250 1686.755 5.265 ;
        RECT 1699.305 5.250 1699.635 5.265 ;
        RECT 1686.425 4.950 1699.635 5.250 ;
        RECT 1686.425 4.935 1686.755 4.950 ;
        RECT 1699.305 4.935 1699.635 4.950 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.850 14.010 1702.990 15.300 ;
        RECT 1702.850 13.870 1703.220 14.010 ;
        RECT 1703.080 5.285 1703.220 13.870 ;
        RECT 1703.010 4.915 1703.290 5.285 ;
        RECT 1716.810 4.915 1717.090 5.285 ;
        RECT 1716.880 2.400 1717.020 4.915 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
      LAYER met3 ;
        RECT 1702.985 5.250 1703.315 5.265 ;
        RECT 1716.785 5.250 1717.115 5.265 ;
        RECT 1702.985 4.950 1717.115 5.250 ;
        RECT 1702.985 4.935 1703.315 4.950 ;
        RECT 1716.785 4.935 1717.115 4.950 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.410 14.010 1719.550 15.300 ;
        RECT 1719.410 13.870 1719.780 14.010 ;
        RECT 1719.640 5.285 1719.780 13.870 ;
        RECT 1719.570 4.915 1719.850 5.285 ;
        RECT 1734.750 4.915 1735.030 5.285 ;
        RECT 1734.820 2.400 1734.960 4.915 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
      LAYER met3 ;
        RECT 1719.545 5.250 1719.875 5.265 ;
        RECT 1734.725 5.250 1735.055 5.265 ;
        RECT 1719.545 4.950 1735.055 5.250 ;
        RECT 1719.545 4.935 1719.875 4.950 ;
        RECT 1734.725 4.935 1735.055 4.950 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.970 14.010 1736.110 15.300 ;
        RECT 1735.970 13.870 1736.340 14.010 ;
        RECT 1736.200 6.645 1736.340 13.870 ;
        RECT 1736.130 6.275 1736.410 6.645 ;
        RECT 1752.230 6.275 1752.510 6.645 ;
        RECT 1752.300 2.400 1752.440 6.275 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
      LAYER met3 ;
        RECT 1736.105 6.610 1736.435 6.625 ;
        RECT 1752.205 6.610 1752.535 6.625 ;
        RECT 1736.105 6.310 1752.535 6.610 ;
        RECT 1736.105 6.295 1736.435 6.310 ;
        RECT 1752.205 6.295 1752.535 6.310 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.530 14.125 1752.670 15.300 ;
        RECT 1752.460 13.755 1752.740 14.125 ;
        RECT 1766.490 13.330 1766.770 13.445 ;
        RECT 1766.490 13.190 1768.080 13.330 ;
        RECT 1766.490 13.075 1766.770 13.190 ;
        RECT 1767.940 1.770 1768.080 13.190 ;
        RECT 1770.030 1.770 1770.590 2.400 ;
        RECT 1767.940 1.630 1770.590 1.770 ;
        RECT 1770.030 -4.800 1770.590 1.630 ;
      LAYER met3 ;
        RECT 1752.435 14.090 1752.765 14.105 ;
        RECT 1752.435 13.790 1762.410 14.090 ;
        RECT 1752.435 13.775 1752.765 13.790 ;
        RECT 1762.110 13.410 1762.410 13.790 ;
        RECT 1766.465 13.410 1766.795 13.425 ;
        RECT 1762.110 13.110 1766.795 13.410 ;
        RECT 1766.465 13.095 1766.795 13.110 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.090 14.805 1769.230 15.300 ;
        RECT 1769.020 14.435 1769.300 14.805 ;
        RECT 1784.430 14.010 1784.710 14.125 ;
        RECT 1784.430 13.870 1785.100 14.010 ;
        RECT 1784.430 13.755 1784.710 13.870 ;
        RECT 1784.960 13.330 1785.100 13.870 ;
        RECT 1784.960 13.190 1787.860 13.330 ;
        RECT 1787.720 2.400 1787.860 13.190 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
      LAYER met3 ;
        RECT 1768.995 14.770 1769.325 14.785 ;
        RECT 1768.995 14.470 1784.490 14.770 ;
        RECT 1768.995 14.455 1769.325 14.470 ;
        RECT 1784.190 14.105 1784.490 14.470 ;
        RECT 1784.190 13.790 1784.735 14.105 ;
        RECT 1784.405 13.775 1784.735 13.790 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1785.650 14.125 1785.790 15.300 ;
        RECT 1785.580 13.755 1785.860 14.125 ;
        RECT 1805.590 13.755 1805.870 14.125 ;
        RECT 1805.660 2.400 1805.800 13.755 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
      LAYER met3 ;
        RECT 1786.950 14.470 1801.050 14.770 ;
        RECT 1785.555 14.090 1785.885 14.105 ;
        RECT 1786.950 14.090 1787.250 14.470 ;
        RECT 1785.555 13.790 1787.250 14.090 ;
        RECT 1800.750 14.090 1801.050 14.470 ;
        RECT 1805.565 14.090 1805.895 14.105 ;
        RECT 1800.750 13.790 1805.895 14.090 ;
        RECT 1785.555 13.775 1785.885 13.790 ;
        RECT 1805.565 13.775 1805.895 13.790 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.210 14.805 1802.350 15.300 ;
        RECT 1802.140 14.435 1802.420 14.805 ;
        RECT 1823.070 13.755 1823.350 14.125 ;
        RECT 1823.140 2.400 1823.280 13.755 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
      LAYER met3 ;
        RECT 1820.950 15.450 1821.330 15.460 ;
        RECT 1817.310 15.150 1821.330 15.450 ;
        RECT 1802.115 14.770 1802.445 14.785 ;
        RECT 1817.310 14.770 1817.610 15.150 ;
        RECT 1820.950 15.140 1821.330 15.150 ;
        RECT 1802.115 14.470 1817.610 14.770 ;
        RECT 1802.115 14.455 1802.445 14.470 ;
        RECT 1820.950 14.090 1821.330 14.100 ;
        RECT 1823.045 14.090 1823.375 14.105 ;
        RECT 1820.950 13.790 1823.375 14.090 ;
        RECT 1820.950 13.780 1821.330 13.790 ;
        RECT 1823.045 13.775 1823.375 13.790 ;
      LAYER met4 ;
        RECT 1820.975 15.135 1821.305 15.465 ;
        RECT 1820.990 14.105 1821.290 15.135 ;
        RECT 1820.975 13.775 1821.305 14.105 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.770 14.805 1818.910 15.300 ;
        RECT 1818.700 14.435 1818.980 14.805 ;
        RECT 1841.010 13.755 1841.290 14.125 ;
        RECT 1841.080 2.400 1841.220 13.755 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
      LAYER met3 ;
        RECT 1818.675 14.770 1819.005 14.785 ;
        RECT 1818.675 14.470 1840.610 14.770 ;
        RECT 1818.675 14.455 1819.005 14.470 ;
        RECT 1840.310 14.090 1840.610 14.470 ;
        RECT 1840.985 14.090 1841.315 14.105 ;
        RECT 1840.310 13.790 1841.315 14.090 ;
        RECT 1840.985 13.775 1841.315 13.790 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1835.240 14.180 1835.560 14.240 ;
        RECT 1856.170 14.180 1856.490 14.240 ;
        RECT 1835.240 14.040 1856.490 14.180 ;
        RECT 1835.240 13.980 1835.560 14.040 ;
        RECT 1856.170 13.980 1856.490 14.040 ;
      LAYER met2 ;
        RECT 1835.330 14.270 1835.470 15.300 ;
        RECT 1835.270 13.950 1835.530 14.270 ;
        RECT 1856.200 13.950 1856.460 14.270 ;
        RECT 1856.260 1.770 1856.400 13.950 ;
        RECT 1858.350 1.770 1858.910 2.400 ;
        RECT 1856.260 1.630 1858.910 1.770 ;
        RECT 1858.350 -4.800 1858.910 1.630 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.050 14.010 792.190 15.300 ;
        RECT 791.820 13.870 792.190 14.010 ;
        RECT 791.820 10.045 791.960 13.870 ;
        RECT 741.610 9.675 741.890 10.045 ;
        RECT 791.750 9.675 792.030 10.045 ;
        RECT 741.680 2.400 741.820 9.675 ;
        RECT 741.470 -4.800 742.030 2.400 ;
      LAYER met3 ;
        RECT 741.585 10.010 741.915 10.025 ;
        RECT 791.725 10.010 792.055 10.025 ;
        RECT 741.585 9.710 792.055 10.010 ;
        RECT 741.585 9.695 741.915 9.710 ;
        RECT 791.725 9.695 792.055 9.710 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1851.800 14.520 1852.120 14.580 ;
        RECT 1875.950 14.520 1876.270 14.580 ;
        RECT 1851.800 14.380 1876.270 14.520 ;
        RECT 1851.800 14.320 1852.120 14.380 ;
        RECT 1875.950 14.320 1876.270 14.380 ;
      LAYER met2 ;
        RECT 1851.890 14.610 1852.030 15.300 ;
        RECT 1851.830 14.290 1852.090 14.610 ;
        RECT 1875.980 14.290 1876.240 14.610 ;
        RECT 1876.040 7.210 1876.180 14.290 ;
        RECT 1876.040 7.070 1876.640 7.210 ;
        RECT 1876.500 2.400 1876.640 7.070 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.450 14.805 1868.590 15.300 ;
        RECT 1868.380 14.435 1868.660 14.805 ;
        RECT 1894.370 13.755 1894.650 14.125 ;
        RECT 1894.440 2.400 1894.580 13.755 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
      LAYER met3 ;
        RECT 1868.355 14.770 1868.685 14.785 ;
        RECT 1868.355 14.470 1893.970 14.770 ;
        RECT 1868.355 14.455 1868.685 14.470 ;
        RECT 1893.670 14.090 1893.970 14.470 ;
        RECT 1894.345 14.090 1894.675 14.105 ;
        RECT 1893.670 13.790 1894.675 14.090 ;
        RECT 1894.345 13.775 1894.675 13.790 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1884.920 14.520 1885.240 14.580 ;
        RECT 1911.370 14.520 1911.690 14.580 ;
        RECT 1884.920 14.380 1911.690 14.520 ;
        RECT 1884.920 14.320 1885.240 14.380 ;
        RECT 1911.370 14.320 1911.690 14.380 ;
      LAYER met2 ;
        RECT 1885.010 14.610 1885.150 15.300 ;
        RECT 1884.950 14.290 1885.210 14.610 ;
        RECT 1911.400 14.290 1911.660 14.610 ;
        RECT 1911.460 7.890 1911.600 14.290 ;
        RECT 1911.460 7.750 1912.060 7.890 ;
        RECT 1911.920 2.400 1912.060 7.750 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1901.710 7.720 1902.030 7.780 ;
        RECT 1928.850 7.720 1929.170 7.780 ;
        RECT 1901.710 7.580 1929.170 7.720 ;
        RECT 1901.710 7.520 1902.030 7.580 ;
        RECT 1928.850 7.520 1929.170 7.580 ;
      LAYER met2 ;
        RECT 1901.570 14.010 1901.710 15.300 ;
        RECT 1901.570 13.870 1901.940 14.010 ;
        RECT 1901.800 7.810 1901.940 13.870 ;
        RECT 1901.740 7.490 1902.000 7.810 ;
        RECT 1928.880 7.490 1929.140 7.810 ;
        RECT 1928.940 3.810 1929.080 7.490 ;
        RECT 1928.940 3.670 1930.000 3.810 ;
        RECT 1929.860 2.400 1930.000 3.670 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.130 14.010 1918.270 15.300 ;
        RECT 1917.900 13.870 1918.270 14.010 ;
        RECT 1917.900 12.765 1918.040 13.870 ;
        RECT 1917.830 12.395 1918.110 12.765 ;
        RECT 1947.270 12.395 1947.550 12.765 ;
        RECT 1947.340 2.400 1947.480 12.395 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER met3 ;
        RECT 1917.550 18.850 1917.930 18.860 ;
        RECT 1946.990 18.850 1947.370 18.860 ;
        RECT 1917.550 18.550 1947.370 18.850 ;
        RECT 1917.550 18.540 1917.930 18.550 ;
        RECT 1946.990 18.540 1947.370 18.550 ;
        RECT 1917.805 12.740 1918.135 12.745 ;
        RECT 1947.245 12.740 1947.575 12.745 ;
        RECT 1917.550 12.730 1918.135 12.740 ;
        RECT 1917.350 12.430 1918.135 12.730 ;
        RECT 1917.550 12.420 1918.135 12.430 ;
        RECT 1946.990 12.730 1947.575 12.740 ;
        RECT 1946.990 12.430 1947.800 12.730 ;
        RECT 1946.990 12.420 1947.575 12.430 ;
        RECT 1917.805 12.415 1918.135 12.420 ;
        RECT 1947.245 12.415 1947.575 12.420 ;
      LAYER met4 ;
        RECT 1917.575 18.535 1917.905 18.865 ;
        RECT 1947.015 18.535 1947.345 18.865 ;
        RECT 1917.590 12.745 1917.890 18.535 ;
        RECT 1947.030 12.745 1947.330 18.535 ;
        RECT 1917.575 12.415 1917.905 12.745 ;
        RECT 1947.015 12.415 1947.345 12.745 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1934.830 7.720 1935.150 7.780 ;
        RECT 1963.350 7.720 1963.670 7.780 ;
        RECT 1934.830 7.580 1963.670 7.720 ;
        RECT 1934.830 7.520 1935.150 7.580 ;
        RECT 1963.350 7.520 1963.670 7.580 ;
      LAYER met2 ;
        RECT 1934.690 14.010 1934.830 15.300 ;
        RECT 1934.690 13.870 1935.060 14.010 ;
        RECT 1934.920 7.810 1935.060 13.870 ;
        RECT 1934.860 7.490 1935.120 7.810 ;
        RECT 1963.380 7.490 1963.640 7.810 ;
        RECT 1963.440 1.770 1963.580 7.490 ;
        RECT 1965.070 1.770 1965.630 2.400 ;
        RECT 1963.440 1.630 1965.630 1.770 ;
        RECT 1965.070 -4.800 1965.630 1.630 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.250 14.010 1951.390 15.300 ;
        RECT 1951.250 13.870 1951.620 14.010 ;
        RECT 1951.480 0.525 1951.620 13.870 ;
        RECT 1951.410 0.155 1951.690 0.525 ;
        RECT 1980.850 0.410 1981.130 0.525 ;
        RECT 1982.550 0.410 1983.110 2.400 ;
        RECT 1980.850 0.270 1983.110 0.410 ;
        RECT 1980.850 0.155 1981.130 0.270 ;
        RECT 1982.550 -4.800 1983.110 0.270 ;
      LAYER met3 ;
        RECT 1951.385 0.490 1951.715 0.505 ;
        RECT 1980.825 0.490 1981.155 0.505 ;
        RECT 1951.385 0.190 1981.155 0.490 ;
        RECT 1951.385 0.175 1951.715 0.190 ;
        RECT 1980.825 0.175 1981.155 0.190 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1967.950 7.720 1968.270 7.780 ;
        RECT 1999.690 7.720 2000.010 7.780 ;
        RECT 1967.950 7.580 2000.010 7.720 ;
        RECT 1967.950 7.520 1968.270 7.580 ;
        RECT 1999.690 7.520 2000.010 7.580 ;
      LAYER met2 ;
        RECT 1967.810 14.690 1967.950 15.300 ;
        RECT 1967.810 14.550 1968.180 14.690 ;
        RECT 1968.040 7.810 1968.180 14.550 ;
        RECT 1967.980 7.490 1968.240 7.810 ;
        RECT 1999.720 7.490 1999.980 7.810 ;
        RECT 1999.780 3.130 1999.920 7.490 ;
        RECT 1999.780 2.990 2000.840 3.130 ;
        RECT 2000.700 2.400 2000.840 2.990 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.370 14.125 1984.510 15.300 ;
        RECT 1984.300 13.755 1984.580 14.125 ;
        RECT 2018.110 13.755 2018.390 14.125 ;
        RECT 2018.180 2.400 2018.320 13.755 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
      LAYER met3 ;
        RECT 1984.275 14.090 1984.605 14.105 ;
        RECT 2018.085 14.090 2018.415 14.105 ;
        RECT 1984.275 13.790 1992.410 14.090 ;
        RECT 1984.275 13.775 1984.605 13.790 ;
        RECT 1992.110 12.730 1992.410 13.790 ;
        RECT 1994.870 13.790 2018.415 14.090 ;
        RECT 1994.870 12.730 1995.170 13.790 ;
        RECT 2018.085 13.775 2018.415 13.790 ;
        RECT 1992.110 12.430 1995.170 12.730 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.930 14.010 2001.070 15.300 ;
        RECT 2000.700 13.870 2001.070 14.010 ;
        RECT 2000.700 4.605 2000.840 13.870 ;
        RECT 2000.630 4.235 2000.910 4.605 ;
        RECT 2036.050 2.875 2036.330 3.245 ;
        RECT 2036.120 2.400 2036.260 2.875 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
      LAYER met3 ;
        RECT 2000.605 4.570 2000.935 4.585 ;
        RECT 2000.605 4.270 2014.950 4.570 ;
        RECT 2000.605 4.255 2000.935 4.270 ;
        RECT 2014.650 3.210 2014.950 4.270 ;
        RECT 2036.025 3.210 2036.355 3.225 ;
        RECT 2014.650 2.910 2036.355 3.210 ;
        RECT 2036.025 2.895 2036.355 2.910 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.610 14.010 808.750 15.300 ;
        RECT 808.380 13.870 808.750 14.010 ;
        RECT 808.380 9.365 808.520 13.870 ;
        RECT 759.090 8.995 759.370 9.365 ;
        RECT 808.310 8.995 808.590 9.365 ;
        RECT 759.160 2.400 759.300 8.995 ;
        RECT 758.950 -4.800 759.510 2.400 ;
      LAYER met3 ;
        RECT 759.065 9.330 759.395 9.345 ;
        RECT 808.285 9.330 808.615 9.345 ;
        RECT 759.065 9.030 808.615 9.330 ;
        RECT 759.065 9.015 759.395 9.030 ;
        RECT 808.285 9.015 808.615 9.030 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.490 14.805 2017.630 15.300 ;
        RECT 2017.420 14.435 2017.700 14.805 ;
        RECT 2052.150 13.330 2052.430 13.445 ;
        RECT 2052.150 13.190 2054.200 13.330 ;
        RECT 2052.150 13.075 2052.430 13.190 ;
        RECT 2054.060 2.400 2054.200 13.190 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
      LAYER met3 ;
        RECT 2017.395 14.770 2017.725 14.785 ;
        RECT 2017.395 14.470 2043.010 14.770 ;
        RECT 2017.395 14.455 2017.725 14.470 ;
        RECT 2042.710 13.410 2043.010 14.470 ;
        RECT 2052.125 13.410 2052.455 13.425 ;
        RECT 2042.710 13.110 2052.455 13.410 ;
        RECT 2052.125 13.095 2052.455 13.110 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.050 14.010 2034.190 15.300 ;
        RECT 2034.050 13.870 2034.420 14.010 ;
        RECT 2034.280 6.645 2034.420 13.870 ;
        RECT 2034.210 6.275 2034.490 6.645 ;
        RECT 2071.470 6.275 2071.750 6.645 ;
        RECT 2071.540 2.400 2071.680 6.275 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
      LAYER met3 ;
        RECT 2034.185 6.610 2034.515 6.625 ;
        RECT 2071.445 6.610 2071.775 6.625 ;
        RECT 2034.185 6.310 2071.775 6.610 ;
        RECT 2034.185 6.295 2034.515 6.310 ;
        RECT 2071.445 6.295 2071.775 6.310 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.610 14.125 2050.750 15.300 ;
        RECT 2050.540 13.755 2050.820 14.125 ;
        RECT 2089.870 13.755 2090.150 14.125 ;
        RECT 2089.940 3.130 2090.080 13.755 ;
        RECT 2089.480 2.990 2090.080 3.130 ;
        RECT 2089.480 2.400 2089.620 2.990 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
      LAYER met3 ;
        RECT 2050.515 14.090 2050.845 14.105 ;
        RECT 2089.845 14.090 2090.175 14.105 ;
        RECT 2050.515 13.790 2073.370 14.090 ;
        RECT 2050.515 13.775 2050.845 13.790 ;
        RECT 2073.070 13.410 2073.370 13.790 ;
        RECT 2084.110 13.790 2090.175 14.090 ;
        RECT 2084.110 13.410 2084.410 13.790 ;
        RECT 2089.845 13.775 2090.175 13.790 ;
        RECT 2073.070 13.110 2084.410 13.410 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.170 14.010 2067.310 15.300 ;
        RECT 2067.170 13.870 2067.540 14.010 ;
        RECT 2067.400 5.285 2067.540 13.870 ;
        RECT 2067.330 4.915 2067.610 5.285 ;
        RECT 2106.890 4.915 2107.170 5.285 ;
        RECT 2106.960 2.400 2107.100 4.915 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
      LAYER met3 ;
        RECT 2067.305 5.250 2067.635 5.265 ;
        RECT 2106.865 5.250 2107.195 5.265 ;
        RECT 2067.305 4.950 2107.195 5.250 ;
        RECT 2067.305 4.935 2067.635 4.950 ;
        RECT 2106.865 4.935 2107.195 4.950 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.730 14.010 2083.870 15.300 ;
        RECT 2083.500 13.870 2083.870 14.010 ;
        RECT 2083.500 5.965 2083.640 13.870 ;
        RECT 2083.430 5.595 2083.710 5.965 ;
        RECT 2124.830 5.595 2125.110 5.965 ;
        RECT 2124.900 2.400 2125.040 5.595 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
      LAYER met3 ;
        RECT 2083.405 5.930 2083.735 5.945 ;
        RECT 2124.805 5.930 2125.135 5.945 ;
        RECT 2083.405 5.630 2125.135 5.930 ;
        RECT 2083.405 5.615 2083.735 5.630 ;
        RECT 2124.805 5.615 2125.135 5.630 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.290 14.010 2100.430 15.300 ;
        RECT 2100.290 13.870 2100.660 14.010 ;
        RECT 2100.520 3.245 2100.660 13.870 ;
        RECT 2100.450 2.875 2100.730 3.245 ;
        RECT 2142.310 2.875 2142.590 3.245 ;
        RECT 2142.380 2.400 2142.520 2.875 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
      LAYER met3 ;
        RECT 2100.425 3.210 2100.755 3.225 ;
        RECT 2142.285 3.210 2142.615 3.225 ;
        RECT 2100.425 2.910 2142.615 3.210 ;
        RECT 2100.425 2.895 2100.755 2.910 ;
        RECT 2142.285 2.895 2142.615 2.910 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2116.850 14.125 2116.990 15.300 ;
        RECT 2116.780 13.755 2117.060 14.125 ;
        RECT 2160.250 13.755 2160.530 14.125 ;
        RECT 2160.320 2.400 2160.460 13.755 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
      LAYER met3 ;
        RECT 2116.755 14.090 2117.085 14.105 ;
        RECT 2160.225 14.090 2160.555 14.105 ;
        RECT 2116.755 13.790 2145.130 14.090 ;
        RECT 2116.755 13.775 2117.085 13.790 ;
        RECT 2144.830 12.730 2145.130 13.790 ;
        RECT 2146.670 13.790 2160.555 14.090 ;
        RECT 2146.670 12.730 2146.970 13.790 ;
        RECT 2160.225 13.775 2160.555 13.790 ;
        RECT 2144.830 12.430 2146.970 12.730 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.410 14.010 2133.550 15.300 ;
        RECT 2133.410 13.870 2133.780 14.010 ;
        RECT 2133.640 1.205 2133.780 13.870 ;
        RECT 2176.880 2.990 2177.940 3.130 ;
        RECT 2176.880 1.205 2177.020 2.990 ;
        RECT 2177.800 2.400 2177.940 2.990 ;
        RECT 2133.570 0.835 2133.850 1.205 ;
        RECT 2176.810 0.835 2177.090 1.205 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
      LAYER met3 ;
        RECT 2133.545 1.170 2133.875 1.185 ;
        RECT 2176.785 1.170 2177.115 1.185 ;
        RECT 2133.545 0.870 2177.115 1.170 ;
        RECT 2133.545 0.855 2133.875 0.870 ;
        RECT 2176.785 0.855 2177.115 0.870 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.970 14.010 2150.110 15.300 ;
        RECT 2149.970 13.870 2150.340 14.010 ;
        RECT 2150.200 12.765 2150.340 13.870 ;
        RECT 2150.130 12.395 2150.410 12.765 ;
        RECT 2195.670 12.395 2195.950 12.765 ;
        RECT 2195.740 2.400 2195.880 12.395 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
      LAYER met3 ;
        RECT 2150.105 12.730 2150.435 12.745 ;
        RECT 2195.645 12.730 2195.975 12.745 ;
        RECT 2150.105 12.430 2195.975 12.730 ;
        RECT 2150.105 12.415 2150.435 12.430 ;
        RECT 2195.645 12.415 2195.975 12.430 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.530 14.010 2166.670 15.300 ;
        RECT 2166.300 13.870 2166.670 14.010 ;
        RECT 2166.300 12.085 2166.440 13.870 ;
        RECT 2166.230 11.715 2166.510 12.085 ;
        RECT 2213.150 11.715 2213.430 12.085 ;
        RECT 2213.220 2.400 2213.360 11.715 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
      LAYER met3 ;
        RECT 2166.205 12.050 2166.535 12.065 ;
        RECT 2213.125 12.050 2213.455 12.065 ;
        RECT 2166.205 11.750 2213.455 12.050 ;
        RECT 2166.205 11.735 2166.535 11.750 ;
        RECT 2213.125 11.735 2213.455 11.750 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.170 14.010 825.310 15.300 ;
        RECT 824.940 13.870 825.310 14.010 ;
        RECT 824.940 11.405 825.080 13.870 ;
        RECT 777.030 11.035 777.310 11.405 ;
        RECT 824.870 11.035 825.150 11.405 ;
        RECT 777.100 2.400 777.240 11.035 ;
        RECT 776.890 -4.800 777.450 2.400 ;
      LAYER met3 ;
        RECT 777.005 11.370 777.335 11.385 ;
        RECT 824.845 11.370 825.175 11.385 ;
        RECT 777.005 11.070 825.175 11.370 ;
        RECT 777.005 11.055 777.335 11.070 ;
        RECT 824.845 11.055 825.175 11.070 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.090 14.010 2183.230 15.300 ;
        RECT 2183.090 13.870 2183.460 14.010 ;
        RECT 2183.320 10.725 2183.460 13.870 ;
        RECT 2183.250 10.355 2183.530 10.725 ;
        RECT 2231.090 10.355 2231.370 10.725 ;
        RECT 2231.160 2.400 2231.300 10.355 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
      LAYER met3 ;
        RECT 2183.225 10.690 2183.555 10.705 ;
        RECT 2231.065 10.690 2231.395 10.705 ;
        RECT 2183.225 10.390 2231.395 10.690 ;
        RECT 2183.225 10.375 2183.555 10.390 ;
        RECT 2231.065 10.375 2231.395 10.390 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.650 14.010 2199.790 15.300 ;
        RECT 2199.650 13.870 2200.020 14.010 ;
        RECT 2199.880 9.365 2200.020 13.870 ;
        RECT 2199.810 8.995 2200.090 9.365 ;
        RECT 2249.030 8.995 2249.310 9.365 ;
        RECT 2249.100 2.400 2249.240 8.995 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
      LAYER met3 ;
        RECT 2199.785 9.330 2200.115 9.345 ;
        RECT 2249.005 9.330 2249.335 9.345 ;
        RECT 2199.785 9.030 2249.335 9.330 ;
        RECT 2199.785 9.015 2200.115 9.030 ;
        RECT 2249.005 9.015 2249.335 9.030 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.210 14.010 2216.350 15.300 ;
        RECT 2216.210 13.870 2216.580 14.010 ;
        RECT 2216.440 12.085 2216.580 13.870 ;
        RECT 2216.370 11.715 2216.650 12.085 ;
        RECT 2266.510 11.715 2266.790 12.085 ;
        RECT 2266.580 2.400 2266.720 11.715 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
      LAYER met3 ;
        RECT 2216.345 12.050 2216.675 12.065 ;
        RECT 2266.485 12.050 2266.815 12.065 ;
        RECT 2216.345 11.750 2266.815 12.050 ;
        RECT 2216.345 11.735 2216.675 11.750 ;
        RECT 2266.485 11.735 2266.815 11.750 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.770 14.010 2232.910 15.300 ;
        RECT 2232.770 13.870 2233.140 14.010 ;
        RECT 2233.000 10.725 2233.140 13.870 ;
        RECT 2232.930 10.355 2233.210 10.725 ;
        RECT 2284.450 10.355 2284.730 10.725 ;
        RECT 2284.520 2.400 2284.660 10.355 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
      LAYER met3 ;
        RECT 2232.905 10.690 2233.235 10.705 ;
        RECT 2284.425 10.690 2284.755 10.705 ;
        RECT 2232.905 10.390 2284.755 10.690 ;
        RECT 2232.905 10.375 2233.235 10.390 ;
        RECT 2284.425 10.375 2284.755 10.390 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2249.240 14.180 2249.560 14.240 ;
        RECT 2301.910 14.180 2302.230 14.240 ;
        RECT 2249.240 14.040 2302.230 14.180 ;
        RECT 2249.240 13.980 2249.560 14.040 ;
        RECT 2301.910 13.980 2302.230 14.040 ;
      LAYER met2 ;
        RECT 2249.330 14.270 2249.470 15.300 ;
        RECT 2249.270 13.950 2249.530 14.270 ;
        RECT 2301.940 13.950 2302.200 14.270 ;
        RECT 2302.000 2.400 2302.140 13.950 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2265.890 14.805 2266.030 15.300 ;
        RECT 2265.820 14.435 2266.100 14.805 ;
        RECT 2319.870 13.755 2320.150 14.125 ;
        RECT 2319.940 2.400 2320.080 13.755 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
      LAYER met3 ;
        RECT 2318.670 17.490 2319.050 17.500 ;
        RECT 2275.470 17.190 2319.050 17.490 ;
        RECT 2265.795 14.770 2266.125 14.785 ;
        RECT 2275.470 14.770 2275.770 17.190 ;
        RECT 2318.670 17.180 2319.050 17.190 ;
        RECT 2265.795 14.470 2275.770 14.770 ;
        RECT 2265.795 14.455 2266.125 14.470 ;
        RECT 2318.670 14.090 2319.050 14.100 ;
        RECT 2319.845 14.090 2320.175 14.105 ;
        RECT 2318.670 13.790 2320.175 14.090 ;
        RECT 2318.670 13.780 2319.050 13.790 ;
        RECT 2319.845 13.775 2320.175 13.790 ;
      LAYER met4 ;
        RECT 2318.695 17.175 2319.025 17.505 ;
        RECT 2318.710 14.105 2319.010 17.175 ;
        RECT 2318.695 13.775 2319.025 14.105 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.450 14.805 2282.590 15.300 ;
        RECT 2282.380 14.435 2282.660 14.805 ;
        RECT 2336.430 12.650 2336.710 12.765 ;
        RECT 2336.430 12.510 2337.560 12.650 ;
        RECT 2336.430 12.395 2336.710 12.510 ;
        RECT 2337.420 2.400 2337.560 12.510 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
      LAYER met3 ;
        RECT 2291.990 16.810 2292.370 16.820 ;
        RECT 2336.150 16.810 2336.530 16.820 ;
        RECT 2291.990 16.510 2336.530 16.810 ;
        RECT 2291.990 16.500 2292.370 16.510 ;
        RECT 2336.150 16.500 2336.530 16.510 ;
        RECT 2282.355 14.770 2282.685 14.785 ;
        RECT 2291.990 14.770 2292.370 14.780 ;
        RECT 2282.355 14.470 2292.370 14.770 ;
        RECT 2282.355 14.455 2282.685 14.470 ;
        RECT 2291.990 14.460 2292.370 14.470 ;
        RECT 2336.405 12.740 2336.735 12.745 ;
        RECT 2336.150 12.730 2336.735 12.740 ;
        RECT 2336.150 12.430 2336.960 12.730 ;
        RECT 2336.150 12.420 2336.735 12.430 ;
        RECT 2336.405 12.415 2336.735 12.420 ;
      LAYER met4 ;
        RECT 2292.015 16.495 2292.345 16.825 ;
        RECT 2336.175 16.495 2336.505 16.825 ;
        RECT 2292.030 14.785 2292.330 16.495 ;
        RECT 2292.015 14.455 2292.345 14.785 ;
        RECT 2336.190 12.745 2336.490 16.495 ;
        RECT 2336.175 12.415 2336.505 12.745 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.010 14.805 2299.150 15.300 ;
        RECT 2298.940 14.435 2299.220 14.805 ;
        RECT 2355.290 13.755 2355.570 14.125 ;
        RECT 2355.360 2.400 2355.500 13.755 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
      LAYER met3 ;
        RECT 2352.750 16.510 2355.810 16.810 ;
        RECT 2352.750 16.130 2353.050 16.510 ;
        RECT 2332.510 15.830 2353.050 16.130 ;
        RECT 2332.510 15.450 2332.810 15.830 ;
        RECT 2319.630 15.150 2332.810 15.450 ;
        RECT 2298.915 14.770 2299.245 14.785 ;
        RECT 2319.630 14.770 2319.930 15.150 ;
        RECT 2298.915 14.470 2319.930 14.770 ;
        RECT 2298.915 14.455 2299.245 14.470 ;
        RECT 2355.510 14.105 2355.810 16.510 ;
        RECT 2355.265 13.790 2355.810 14.105 ;
        RECT 2355.265 13.775 2355.595 13.790 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.570 13.870 2315.710 15.300 ;
        RECT 2315.570 13.730 2315.940 13.870 ;
        RECT 2315.800 11.405 2315.940 13.730 ;
        RECT 2315.730 11.035 2316.010 11.405 ;
        RECT 2372.770 11.035 2373.050 11.405 ;
        RECT 2372.840 2.400 2372.980 11.035 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
      LAYER met3 ;
        RECT 2315.705 11.370 2316.035 11.385 ;
        RECT 2372.745 11.370 2373.075 11.385 ;
        RECT 2315.705 11.070 2373.075 11.370 ;
        RECT 2315.705 11.055 2316.035 11.070 ;
        RECT 2372.745 11.055 2373.075 11.070 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2331.810 6.020 2332.130 6.080 ;
        RECT 2389.310 6.020 2389.630 6.080 ;
        RECT 2331.810 5.880 2389.630 6.020 ;
        RECT 2331.810 5.820 2332.130 5.880 ;
        RECT 2389.310 5.820 2389.630 5.880 ;
      LAYER met2 ;
        RECT 2332.130 13.870 2332.270 15.300 ;
        RECT 2331.900 13.730 2332.270 13.870 ;
        RECT 2331.900 6.110 2332.040 13.730 ;
        RECT 2331.840 5.790 2332.100 6.110 ;
        RECT 2389.340 5.790 2389.600 6.110 ;
        RECT 2389.400 3.130 2389.540 5.790 ;
        RECT 2389.400 2.990 2390.920 3.130 ;
        RECT 2390.780 2.400 2390.920 2.990 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.730 14.010 841.870 15.300 ;
        RECT 840.120 13.870 841.870 14.010 ;
        RECT 794.370 0.410 794.930 2.400 ;
        RECT 840.120 0.525 840.260 13.870 ;
        RECT 796.350 0.410 796.630 0.525 ;
        RECT 794.370 0.270 796.630 0.410 ;
        RECT 794.370 -4.800 794.930 0.270 ;
        RECT 796.350 0.155 796.630 0.270 ;
        RECT 840.050 0.155 840.330 0.525 ;
      LAYER met3 ;
        RECT 796.325 0.490 796.655 0.505 ;
        RECT 840.025 0.490 840.355 0.505 ;
        RECT 796.325 0.190 840.355 0.490 ;
        RECT 796.325 0.175 796.655 0.190 ;
        RECT 840.025 0.175 840.355 0.190 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 0.920 642.090 0.980 ;
        RECT 697.890 0.920 698.210 0.980 ;
        RECT 641.770 0.780 698.210 0.920 ;
        RECT 641.770 0.720 642.090 0.780 ;
        RECT 697.890 0.720 698.210 0.780 ;
      LAYER met2 ;
        RECT 698.210 14.010 698.350 15.300 ;
        RECT 697.980 13.870 698.350 14.010 ;
        RECT 640.730 1.090 641.290 2.400 ;
        RECT 640.730 1.010 642.000 1.090 ;
        RECT 697.980 1.010 698.120 13.870 ;
        RECT 640.730 0.950 642.060 1.010 ;
        RECT 640.730 -4.800 641.290 0.950 ;
        RECT 641.800 0.690 642.060 0.950 ;
        RECT 697.920 0.690 698.180 1.010 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2354.210 14.690 2354.350 15.300 ;
        RECT 2354.210 14.550 2356.420 14.690 ;
        RECT 2356.280 14.125 2356.420 14.550 ;
        RECT 2356.210 13.755 2356.490 14.125 ;
        RECT 2414.170 13.755 2414.450 14.125 ;
        RECT 2414.240 2.400 2414.380 13.755 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
      LAYER met3 ;
        RECT 2356.185 14.090 2356.515 14.105 ;
        RECT 2414.145 14.090 2414.475 14.105 ;
        RECT 2356.185 13.790 2414.475 14.090 ;
        RECT 2356.185 13.775 2356.515 13.790 ;
        RECT 2414.145 13.775 2414.475 13.790 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2370.910 0.920 2371.230 0.980 ;
        RECT 2433.010 0.920 2433.330 0.980 ;
        RECT 2370.910 0.780 2433.330 0.920 ;
        RECT 2370.910 0.720 2371.230 0.780 ;
        RECT 2433.010 0.720 2433.330 0.780 ;
      LAYER met2 ;
        RECT 2370.770 14.010 2370.910 15.300 ;
        RECT 2370.770 13.870 2371.140 14.010 ;
        RECT 2371.000 1.010 2371.140 13.870 ;
        RECT 2431.970 1.090 2432.530 2.400 ;
        RECT 2431.970 1.010 2433.240 1.090 ;
        RECT 2370.940 0.690 2371.200 1.010 ;
        RECT 2431.970 0.950 2433.300 1.010 ;
        RECT 2431.970 -4.800 2432.530 0.950 ;
        RECT 2433.040 0.690 2433.300 0.950 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2387.010 0.580 2387.330 0.640 ;
        RECT 2450.490 0.580 2450.810 0.640 ;
        RECT 2387.010 0.440 2450.810 0.580 ;
        RECT 2387.010 0.380 2387.330 0.440 ;
        RECT 2450.490 0.380 2450.810 0.440 ;
      LAYER met2 ;
        RECT 2387.330 14.010 2387.470 15.300 ;
        RECT 2387.100 13.870 2387.470 14.010 ;
        RECT 2387.100 0.670 2387.240 13.870 ;
        RECT 2387.040 0.350 2387.300 0.670 ;
        RECT 2449.450 0.410 2450.010 2.400 ;
        RECT 2450.520 0.410 2450.780 0.670 ;
        RECT 2449.450 0.350 2450.780 0.410 ;
        RECT 2449.450 0.270 2450.720 0.350 ;
        RECT 2449.450 -4.800 2450.010 0.270 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2403.890 14.010 2404.030 15.300 ;
        RECT 2403.890 13.870 2404.260 14.010 ;
        RECT 2404.120 3.245 2404.260 13.870 ;
        RECT 2404.050 2.875 2404.330 3.245 ;
        RECT 2467.530 2.875 2467.810 3.245 ;
        RECT 2467.600 2.400 2467.740 2.875 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
      LAYER met3 ;
        RECT 2404.025 3.210 2404.355 3.225 ;
        RECT 2467.505 3.210 2467.835 3.225 ;
        RECT 2404.025 2.910 2467.835 3.210 ;
        RECT 2404.025 2.895 2404.355 2.910 ;
        RECT 2467.505 2.895 2467.835 2.910 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2421.050 1.260 2421.370 1.320 ;
        RECT 2486.370 1.260 2486.690 1.320 ;
        RECT 2421.050 1.120 2486.690 1.260 ;
        RECT 2421.050 1.060 2421.370 1.120 ;
        RECT 2486.370 1.060 2486.690 1.120 ;
      LAYER met2 ;
        RECT 2420.450 14.010 2420.590 15.300 ;
        RECT 2420.450 13.870 2421.280 14.010 ;
        RECT 2421.140 1.350 2421.280 13.870 ;
        RECT 2421.080 1.030 2421.340 1.350 ;
        RECT 2485.330 1.090 2485.890 2.400 ;
        RECT 2486.400 1.090 2486.660 1.350 ;
        RECT 2485.330 1.030 2486.660 1.090 ;
        RECT 2485.330 0.950 2486.600 1.030 ;
        RECT 2485.330 -4.800 2485.890 0.950 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.010 14.010 2437.150 15.300 ;
        RECT 2436.320 13.870 2437.150 14.010 ;
        RECT 2436.320 1.205 2436.460 13.870 ;
        RECT 2501.640 2.990 2503.160 3.130 ;
        RECT 2501.640 1.205 2501.780 2.990 ;
        RECT 2503.020 2.400 2503.160 2.990 ;
        RECT 2436.250 0.835 2436.530 1.205 ;
        RECT 2501.570 0.835 2501.850 1.205 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
      LAYER met3 ;
        RECT 2436.225 1.170 2436.555 1.185 ;
        RECT 2501.545 1.170 2501.875 1.185 ;
        RECT 2436.225 0.870 2501.875 1.170 ;
        RECT 2436.225 0.855 2436.555 0.870 ;
        RECT 2501.545 0.855 2501.875 0.870 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2453.250 0.920 2453.570 0.980 ;
        RECT 2519.030 0.920 2519.350 0.980 ;
        RECT 2453.250 0.780 2519.350 0.920 ;
        RECT 2453.250 0.720 2453.570 0.780 ;
        RECT 2519.030 0.720 2519.350 0.780 ;
      LAYER met2 ;
        RECT 2453.570 14.010 2453.710 15.300 ;
        RECT 2453.340 13.870 2453.710 14.010 ;
        RECT 2453.340 1.010 2453.480 13.870 ;
        RECT 2520.750 1.090 2521.310 2.400 ;
        RECT 2519.120 1.010 2521.310 1.090 ;
        RECT 2453.280 0.690 2453.540 1.010 ;
        RECT 2519.060 0.950 2521.310 1.010 ;
        RECT 2519.060 0.690 2519.320 0.950 ;
        RECT 2520.750 -4.800 2521.310 0.950 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2469.810 0.580 2470.130 0.640 ;
        RECT 2536.510 0.580 2536.830 0.640 ;
        RECT 2469.810 0.440 2536.830 0.580 ;
        RECT 2469.810 0.380 2470.130 0.440 ;
        RECT 2536.510 0.380 2536.830 0.440 ;
      LAYER met2 ;
        RECT 2470.130 14.010 2470.270 15.300 ;
        RECT 2469.900 13.870 2470.270 14.010 ;
        RECT 2469.900 0.670 2470.040 13.870 ;
        RECT 2469.840 0.350 2470.100 0.670 ;
        RECT 2536.540 0.410 2536.800 0.670 ;
        RECT 2538.230 0.410 2538.790 2.400 ;
        RECT 2536.540 0.350 2538.790 0.410 ;
        RECT 2536.600 0.270 2538.790 0.350 ;
        RECT 2538.230 -4.800 2538.790 0.270 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2486.830 3.640 2487.150 3.700 ;
        RECT 2486.830 3.500 2522.020 3.640 ;
        RECT 2486.830 3.440 2487.150 3.500 ;
        RECT 2521.880 2.280 2522.020 3.500 ;
        RECT 2557.210 2.280 2557.530 2.340 ;
        RECT 2521.880 2.140 2557.530 2.280 ;
        RECT 2557.210 2.080 2557.530 2.140 ;
      LAYER met2 ;
        RECT 2486.690 14.010 2486.830 15.300 ;
        RECT 2486.690 13.870 2487.060 14.010 ;
        RECT 2486.920 3.730 2487.060 13.870 ;
        RECT 2486.860 3.410 2487.120 3.730 ;
        RECT 2556.170 1.770 2556.730 2.400 ;
        RECT 2557.240 2.050 2557.500 2.370 ;
        RECT 2557.300 1.770 2557.440 2.050 ;
        RECT 2556.170 1.630 2557.440 1.770 ;
        RECT 2556.170 -4.800 2556.730 1.630 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2503.390 3.980 2503.710 4.040 ;
        RECT 2573.770 3.980 2574.090 4.040 ;
        RECT 2503.390 3.840 2574.090 3.980 ;
        RECT 2503.390 3.780 2503.710 3.840 ;
        RECT 2573.770 3.780 2574.090 3.840 ;
      LAYER met2 ;
        RECT 2503.250 14.010 2503.390 15.300 ;
        RECT 2503.250 13.870 2503.620 14.010 ;
        RECT 2503.480 4.070 2503.620 13.870 ;
        RECT 2503.420 3.750 2503.680 4.070 ;
        RECT 2573.800 3.750 2574.060 4.070 ;
        RECT 2573.860 2.400 2574.000 3.750 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 820.710 6.700 821.030 6.760 ;
        RECT 863.490 6.700 863.810 6.760 ;
        RECT 820.710 6.560 863.810 6.700 ;
        RECT 820.710 6.500 821.030 6.560 ;
        RECT 863.490 6.500 863.810 6.560 ;
      LAYER met2 ;
        RECT 863.810 14.010 863.950 15.300 ;
        RECT 863.580 13.870 863.950 14.010 ;
        RECT 863.580 6.790 863.720 13.870 ;
        RECT 820.740 6.470 821.000 6.790 ;
        RECT 863.520 6.470 863.780 6.790 ;
        RECT 818.290 1.770 818.850 2.400 ;
        RECT 820.800 1.770 820.940 6.470 ;
        RECT 818.290 1.630 820.940 1.770 ;
        RECT 818.290 -4.800 818.850 1.630 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.810 14.010 2519.950 15.300 ;
        RECT 2518.660 13.870 2519.950 14.010 ;
        RECT 2518.660 0.525 2518.800 13.870 ;
        RECT 2590.880 2.990 2591.940 3.130 ;
        RECT 2590.880 0.525 2591.020 2.990 ;
        RECT 2591.800 2.400 2591.940 2.990 ;
        RECT 2518.590 0.155 2518.870 0.525 ;
        RECT 2590.810 0.155 2591.090 0.525 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
      LAYER met3 ;
        RECT 2518.565 0.490 2518.895 0.505 ;
        RECT 2590.785 0.490 2591.115 0.505 ;
        RECT 2518.565 0.190 2591.115 0.490 ;
        RECT 2518.565 0.175 2518.895 0.190 ;
        RECT 2590.785 0.175 2591.115 0.190 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2536.050 0.920 2536.370 0.980 ;
        RECT 2608.270 0.920 2608.590 0.980 ;
        RECT 2536.050 0.780 2608.590 0.920 ;
        RECT 2536.050 0.720 2536.370 0.780 ;
        RECT 2608.270 0.720 2608.590 0.780 ;
      LAYER met2 ;
        RECT 2536.370 14.010 2536.510 15.300 ;
        RECT 2536.140 13.870 2536.510 14.010 ;
        RECT 2536.140 1.010 2536.280 13.870 ;
        RECT 2609.070 1.090 2609.630 2.400 ;
        RECT 2608.360 1.010 2609.630 1.090 ;
        RECT 2536.080 0.690 2536.340 1.010 ;
        RECT 2608.300 0.950 2609.630 1.010 ;
        RECT 2608.300 0.690 2608.560 0.950 ;
        RECT 2609.070 -4.800 2609.630 0.950 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2552.610 0.580 2552.930 0.640 ;
        RECT 2628.050 0.580 2628.370 0.640 ;
        RECT 2552.610 0.440 2628.370 0.580 ;
        RECT 2552.610 0.380 2552.930 0.440 ;
        RECT 2628.050 0.380 2628.370 0.440 ;
      LAYER met2 ;
        RECT 2552.930 14.010 2553.070 15.300 ;
        RECT 2552.700 13.870 2553.070 14.010 ;
        RECT 2552.700 0.670 2552.840 13.870 ;
        RECT 2552.640 0.350 2552.900 0.670 ;
        RECT 2627.010 0.410 2627.570 2.400 ;
        RECT 2628.080 0.410 2628.340 0.670 ;
        RECT 2627.010 0.350 2628.340 0.410 ;
        RECT 2627.010 0.270 2628.280 0.350 ;
        RECT 2627.010 -4.800 2627.570 0.270 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2569.630 3.640 2569.950 3.700 ;
        RECT 2645.070 3.640 2645.390 3.700 ;
        RECT 2569.630 3.500 2645.390 3.640 ;
        RECT 2569.630 3.440 2569.950 3.500 ;
        RECT 2645.070 3.440 2645.390 3.500 ;
      LAYER met2 ;
        RECT 2569.490 14.010 2569.630 15.300 ;
        RECT 2569.490 13.870 2569.860 14.010 ;
        RECT 2569.720 3.730 2569.860 13.870 ;
        RECT 2569.660 3.410 2569.920 3.730 ;
        RECT 2645.100 3.410 2645.360 3.730 ;
        RECT 2645.160 2.400 2645.300 3.410 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2586.650 1.600 2586.970 1.660 ;
        RECT 2660.710 1.600 2661.030 1.660 ;
        RECT 2586.650 1.460 2661.030 1.600 ;
        RECT 2586.650 1.400 2586.970 1.460 ;
        RECT 2660.710 1.400 2661.030 1.460 ;
      LAYER met2 ;
        RECT 2586.050 14.010 2586.190 15.300 ;
        RECT 2586.050 13.870 2586.880 14.010 ;
        RECT 2586.740 1.690 2586.880 13.870 ;
        RECT 2662.430 1.770 2662.990 2.400 ;
        RECT 2660.800 1.690 2662.990 1.770 ;
        RECT 2586.680 1.370 2586.940 1.690 ;
        RECT 2660.740 1.630 2662.990 1.690 ;
        RECT 2660.740 1.370 2661.000 1.630 ;
        RECT 2662.430 -4.800 2662.990 1.630 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2602.750 1.260 2603.070 1.320 ;
        RECT 2681.410 1.260 2681.730 1.320 ;
        RECT 2602.750 1.120 2681.730 1.260 ;
        RECT 2602.750 1.060 2603.070 1.120 ;
        RECT 2681.410 1.060 2681.730 1.120 ;
      LAYER met2 ;
        RECT 2602.610 14.010 2602.750 15.300 ;
        RECT 2602.610 13.870 2602.980 14.010 ;
        RECT 2602.840 1.350 2602.980 13.870 ;
        RECT 2602.780 1.030 2603.040 1.350 ;
        RECT 2680.370 1.090 2680.930 2.400 ;
        RECT 2681.440 1.090 2681.700 1.350 ;
        RECT 2680.370 1.030 2681.700 1.090 ;
        RECT 2680.370 0.950 2681.640 1.030 ;
        RECT 2680.370 -4.800 2680.930 0.950 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2619.310 1.940 2619.630 2.000 ;
        RECT 2698.890 1.940 2699.210 2.000 ;
        RECT 2619.310 1.800 2699.210 1.940 ;
        RECT 2619.310 1.740 2619.630 1.800 ;
        RECT 2698.890 1.740 2699.210 1.800 ;
      LAYER met2 ;
        RECT 2619.170 14.010 2619.310 15.300 ;
        RECT 2619.170 13.870 2619.540 14.010 ;
        RECT 2619.400 2.030 2619.540 13.870 ;
        RECT 2619.340 1.710 2619.600 2.030 ;
        RECT 2697.850 1.770 2698.410 2.400 ;
        RECT 2698.920 1.770 2699.180 2.030 ;
        RECT 2697.850 1.710 2699.180 1.770 ;
        RECT 2697.850 1.630 2699.120 1.710 ;
        RECT 2697.850 -4.800 2698.410 1.630 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2635.410 0.580 2635.730 0.640 ;
        RECT 2714.070 0.580 2714.390 0.640 ;
        RECT 2635.410 0.440 2714.390 0.580 ;
        RECT 2635.410 0.380 2635.730 0.440 ;
        RECT 2714.070 0.380 2714.390 0.440 ;
      LAYER met2 ;
        RECT 2635.730 13.870 2635.870 15.300 ;
        RECT 2635.500 13.730 2635.870 13.870 ;
        RECT 2635.500 0.670 2635.640 13.730 ;
        RECT 2635.440 0.350 2635.700 0.670 ;
        RECT 2714.100 0.410 2714.360 0.670 ;
        RECT 2715.790 0.410 2716.350 2.400 ;
        RECT 2714.100 0.350 2716.350 0.410 ;
        RECT 2714.160 0.270 2716.350 0.350 ;
        RECT 2715.790 -4.800 2716.350 0.270 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2652.430 6.020 2652.750 6.080 ;
        RECT 2732.470 6.020 2732.790 6.080 ;
        RECT 2652.430 5.880 2732.790 6.020 ;
        RECT 2652.430 5.820 2652.750 5.880 ;
        RECT 2732.470 5.820 2732.790 5.880 ;
      LAYER met2 ;
        RECT 2652.290 13.870 2652.430 15.300 ;
        RECT 2652.290 13.730 2652.660 13.870 ;
        RECT 2652.520 6.110 2652.660 13.730 ;
        RECT 2652.460 5.790 2652.720 6.110 ;
        RECT 2732.500 5.790 2732.760 6.110 ;
        RECT 2732.560 1.770 2732.700 5.790 ;
        RECT 2733.270 1.770 2733.830 2.400 ;
        RECT 2732.560 1.630 2733.830 1.770 ;
        RECT 2733.270 -4.800 2733.830 1.630 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2668.990 6.700 2669.310 6.760 ;
        RECT 2750.410 6.700 2750.730 6.760 ;
        RECT 2668.990 6.560 2750.730 6.700 ;
        RECT 2668.990 6.500 2669.310 6.560 ;
        RECT 2750.410 6.500 2750.730 6.560 ;
      LAYER met2 ;
        RECT 2668.850 13.870 2668.990 15.300 ;
        RECT 2668.850 13.730 2669.220 13.870 ;
        RECT 2669.080 6.790 2669.220 13.730 ;
        RECT 2669.020 6.470 2669.280 6.790 ;
        RECT 2750.440 6.470 2750.700 6.790 ;
        RECT 2750.500 3.810 2750.640 6.470 ;
        RECT 2750.500 3.670 2751.560 3.810 ;
        RECT 2751.420 2.400 2751.560 3.670 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.370 14.010 880.510 15.300 ;
        RECT 880.140 13.870 880.510 14.010 ;
        RECT 880.140 3.925 880.280 13.870 ;
        RECT 835.910 3.555 836.190 3.925 ;
        RECT 880.070 3.555 880.350 3.925 ;
        RECT 835.980 2.400 836.120 3.555 ;
        RECT 835.770 -4.800 836.330 2.400 ;
      LAYER met3 ;
        RECT 835.885 3.890 836.215 3.905 ;
        RECT 880.045 3.890 880.375 3.905 ;
        RECT 835.885 3.590 880.375 3.890 ;
        RECT 835.885 3.575 836.215 3.590 ;
        RECT 880.045 3.575 880.375 3.590 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2685.550 6.360 2685.870 6.420 ;
        RECT 2685.550 6.220 2739.370 6.360 ;
        RECT 2685.550 6.160 2685.870 6.220 ;
        RECT 2739.230 6.020 2739.370 6.220 ;
        RECT 2768.810 6.020 2769.130 6.080 ;
        RECT 2739.230 5.880 2769.130 6.020 ;
        RECT 2768.810 5.820 2769.130 5.880 ;
      LAYER met2 ;
        RECT 2685.410 14.010 2685.550 15.300 ;
        RECT 2685.410 13.870 2685.780 14.010 ;
        RECT 2685.640 6.450 2685.780 13.870 ;
        RECT 2685.580 6.130 2685.840 6.450 ;
        RECT 2768.840 5.790 2769.100 6.110 ;
        RECT 2768.900 2.400 2769.040 5.790 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2702.110 0.920 2702.430 0.980 ;
        RECT 2784.910 0.920 2785.230 0.980 ;
        RECT 2702.110 0.780 2785.230 0.920 ;
        RECT 2702.110 0.720 2702.430 0.780 ;
        RECT 2784.910 0.720 2785.230 0.780 ;
      LAYER met2 ;
        RECT 2701.970 14.010 2702.110 15.300 ;
        RECT 2701.970 13.870 2702.340 14.010 ;
        RECT 2702.200 1.010 2702.340 13.870 ;
        RECT 2786.630 1.090 2787.190 2.400 ;
        RECT 2785.000 1.010 2787.190 1.090 ;
        RECT 2702.140 0.690 2702.400 1.010 ;
        RECT 2784.940 0.950 2787.190 1.010 ;
        RECT 2784.940 0.690 2785.200 0.950 ;
        RECT 2786.630 -4.800 2787.190 0.950 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2718.210 0.580 2718.530 0.640 ;
        RECT 2802.390 0.580 2802.710 0.640 ;
        RECT 2718.210 0.440 2802.710 0.580 ;
        RECT 2718.210 0.380 2718.530 0.440 ;
        RECT 2802.390 0.380 2802.710 0.440 ;
      LAYER met2 ;
        RECT 2718.530 14.010 2718.670 15.300 ;
        RECT 2718.300 13.870 2718.670 14.010 ;
        RECT 2718.300 0.670 2718.440 13.870 ;
        RECT 2718.240 0.350 2718.500 0.670 ;
        RECT 2802.420 0.410 2802.680 0.670 ;
        RECT 2804.110 0.410 2804.670 2.400 ;
        RECT 2802.420 0.350 2804.670 0.410 ;
        RECT 2802.480 0.270 2804.670 0.350 ;
        RECT 2804.110 -4.800 2804.670 0.270 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2735.230 1.940 2735.550 2.000 ;
        RECT 2823.090 1.940 2823.410 2.000 ;
        RECT 2735.230 1.800 2823.410 1.940 ;
        RECT 2735.230 1.740 2735.550 1.800 ;
        RECT 2823.090 1.740 2823.410 1.800 ;
      LAYER met2 ;
        RECT 2735.090 13.870 2735.230 15.300 ;
        RECT 2735.090 13.730 2735.460 13.870 ;
        RECT 2735.320 2.030 2735.460 13.730 ;
        RECT 2735.260 1.710 2735.520 2.030 ;
        RECT 2822.050 1.770 2822.610 2.400 ;
        RECT 2823.120 1.770 2823.380 2.030 ;
        RECT 2822.050 1.710 2823.380 1.770 ;
        RECT 2822.050 1.630 2823.320 1.710 ;
        RECT 2822.050 -4.800 2822.610 1.630 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2751.790 6.360 2752.110 6.420 ;
        RECT 2837.810 6.360 2838.130 6.420 ;
        RECT 2751.790 6.220 2838.130 6.360 ;
        RECT 2751.790 6.160 2752.110 6.220 ;
        RECT 2837.810 6.160 2838.130 6.220 ;
      LAYER met2 ;
        RECT 2751.650 13.870 2751.790 15.300 ;
        RECT 2751.650 13.730 2752.020 13.870 ;
        RECT 2751.880 6.450 2752.020 13.730 ;
        RECT 2751.820 6.130 2752.080 6.450 ;
        RECT 2837.840 6.130 2838.100 6.450 ;
        RECT 2837.900 1.770 2838.040 6.130 ;
        RECT 2839.990 1.770 2840.550 2.400 ;
        RECT 2837.900 1.630 2840.550 1.770 ;
        RECT 2839.990 -4.800 2840.550 1.630 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2768.350 6.700 2768.670 6.760 ;
        RECT 2855.290 6.700 2855.610 6.760 ;
        RECT 2768.350 6.560 2855.610 6.700 ;
        RECT 2768.350 6.500 2768.670 6.560 ;
        RECT 2855.290 6.500 2855.610 6.560 ;
      LAYER met2 ;
        RECT 2768.210 14.010 2768.350 15.300 ;
        RECT 2768.210 13.870 2768.580 14.010 ;
        RECT 2768.440 6.790 2768.580 13.870 ;
        RECT 2768.380 6.470 2768.640 6.790 ;
        RECT 2855.320 6.470 2855.580 6.790 ;
        RECT 2855.380 1.770 2855.520 6.470 ;
        RECT 2857.470 1.770 2858.030 2.400 ;
        RECT 2855.380 1.630 2858.030 1.770 ;
        RECT 2857.470 -4.800 2858.030 1.630 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2784.450 1.260 2784.770 1.320 ;
        RECT 2876.450 1.260 2876.770 1.320 ;
        RECT 2784.450 1.120 2876.770 1.260 ;
        RECT 2784.450 1.060 2784.770 1.120 ;
        RECT 2876.450 1.060 2876.770 1.120 ;
      LAYER met2 ;
        RECT 2784.770 14.010 2784.910 15.300 ;
        RECT 2784.540 13.870 2784.910 14.010 ;
        RECT 2784.540 1.350 2784.680 13.870 ;
        RECT 2784.480 1.030 2784.740 1.350 ;
        RECT 2875.410 1.090 2875.970 2.400 ;
        RECT 2876.480 1.090 2876.740 1.350 ;
        RECT 2875.410 1.030 2876.740 1.090 ;
        RECT 2875.410 0.950 2876.680 1.030 ;
        RECT 2875.410 -4.800 2875.970 0.950 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2801.010 0.920 2801.330 0.980 ;
        RECT 2893.930 0.920 2894.250 0.980 ;
        RECT 2801.010 0.780 2894.250 0.920 ;
        RECT 2801.010 0.720 2801.330 0.780 ;
        RECT 2893.930 0.720 2894.250 0.780 ;
      LAYER met2 ;
        RECT 2801.330 14.010 2801.470 15.300 ;
        RECT 2801.100 13.870 2801.470 14.010 ;
        RECT 2801.100 1.010 2801.240 13.870 ;
        RECT 2892.890 1.090 2893.450 2.400 ;
        RECT 2892.890 1.010 2894.160 1.090 ;
        RECT 2801.040 0.690 2801.300 1.010 ;
        RECT 2892.890 0.950 2894.220 1.010 ;
        RECT 2892.890 -4.800 2893.450 0.950 ;
        RECT 2893.960 0.690 2894.220 0.950 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.930 14.010 897.070 15.300 ;
        RECT 896.700 13.870 897.070 14.010 ;
        RECT 896.700 2.565 896.840 13.870 ;
        RECT 852.930 2.195 853.210 2.565 ;
        RECT 853.000 1.770 853.140 2.195 ;
        RECT 853.710 1.770 854.270 2.400 ;
        RECT 896.630 2.195 896.910 2.565 ;
        RECT 853.000 1.630 854.270 1.770 ;
        RECT 853.710 -4.800 854.270 1.630 ;
      LAYER met3 ;
        RECT 852.905 2.530 853.235 2.545 ;
        RECT 896.605 2.530 896.935 2.545 ;
        RECT 852.905 2.230 896.935 2.530 ;
        RECT 852.905 2.215 853.235 2.230 ;
        RECT 896.605 2.215 896.935 2.230 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.490 14.010 913.630 15.300 ;
        RECT 913.260 13.870 913.630 14.010 ;
        RECT 913.260 6.645 913.400 13.870 ;
        RECT 871.330 6.275 871.610 6.645 ;
        RECT 913.190 6.275 913.470 6.645 ;
        RECT 871.400 2.400 871.540 6.275 ;
        RECT 871.190 -4.800 871.750 2.400 ;
      LAYER met3 ;
        RECT 871.305 6.610 871.635 6.625 ;
        RECT 913.165 6.610 913.495 6.625 ;
        RECT 871.305 6.310 913.495 6.610 ;
        RECT 871.305 6.295 871.635 6.310 ;
        RECT 913.165 6.295 913.495 6.310 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.050 14.010 930.190 15.300 ;
        RECT 929.820 13.870 930.190 14.010 ;
        RECT 929.820 5.285 929.960 13.870 ;
        RECT 889.270 4.915 889.550 5.285 ;
        RECT 929.750 4.915 930.030 5.285 ;
        RECT 889.340 2.400 889.480 4.915 ;
        RECT 889.130 -4.800 889.690 2.400 ;
      LAYER met3 ;
        RECT 889.245 5.250 889.575 5.265 ;
        RECT 929.725 5.250 930.055 5.265 ;
        RECT 889.245 4.950 930.055 5.250 ;
        RECT 889.245 4.935 889.575 4.950 ;
        RECT 929.725 4.935 930.055 4.950 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.610 14.010 946.750 15.300 ;
        RECT 946.380 13.870 946.750 14.010 ;
        RECT 946.380 4.605 946.520 13.870 ;
        RECT 907.210 4.235 907.490 4.605 ;
        RECT 946.310 4.235 946.590 4.605 ;
        RECT 907.280 2.400 907.420 4.235 ;
        RECT 907.070 -4.800 907.630 2.400 ;
      LAYER met3 ;
        RECT 907.185 4.570 907.515 4.585 ;
        RECT 946.285 4.570 946.615 4.585 ;
        RECT 907.185 4.270 946.615 4.570 ;
        RECT 907.185 4.255 907.515 4.270 ;
        RECT 946.285 4.255 946.615 4.270 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.170 14.010 963.310 15.300 ;
        RECT 962.940 13.870 963.310 14.010 ;
        RECT 962.940 6.645 963.080 13.870 ;
        RECT 924.690 6.275 924.970 6.645 ;
        RECT 962.870 6.275 963.150 6.645 ;
        RECT 924.760 2.400 924.900 6.275 ;
        RECT 924.550 -4.800 925.110 2.400 ;
      LAYER met3 ;
        RECT 924.665 6.610 924.995 6.625 ;
        RECT 962.845 6.610 963.175 6.625 ;
        RECT 924.665 6.310 963.175 6.610 ;
        RECT 924.665 6.295 924.995 6.310 ;
        RECT 962.845 6.295 963.175 6.310 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.730 14.010 979.870 15.300 ;
        RECT 979.500 13.870 979.870 14.010 ;
        RECT 979.500 3.245 979.640 13.870 ;
        RECT 979.430 2.875 979.710 3.245 ;
        RECT 942.490 1.770 943.050 2.400 ;
        RECT 944.930 1.770 945.210 1.885 ;
        RECT 942.490 1.630 945.210 1.770 ;
        RECT 942.490 -4.800 943.050 1.630 ;
        RECT 944.930 1.515 945.210 1.630 ;
      LAYER met3 ;
        RECT 979.405 3.210 979.735 3.225 ;
        RECT 963.550 2.910 979.735 3.210 ;
        RECT 944.905 1.850 945.235 1.865 ;
        RECT 963.550 1.850 963.850 2.910 ;
        RECT 979.405 2.895 979.735 2.910 ;
        RECT 944.905 1.550 963.850 1.850 ;
        RECT 944.905 1.535 945.235 1.550 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.290 14.010 996.430 15.300 ;
        RECT 996.060 13.870 996.430 14.010 ;
        RECT 996.060 4.605 996.200 13.870 ;
        RECT 960.110 4.235 960.390 4.605 ;
        RECT 995.990 4.235 996.270 4.605 ;
        RECT 960.180 2.400 960.320 4.235 ;
        RECT 959.970 -4.800 960.530 2.400 ;
      LAYER met3 ;
        RECT 960.085 4.570 960.415 4.585 ;
        RECT 995.965 4.570 996.295 4.585 ;
        RECT 960.085 4.270 996.295 4.570 ;
        RECT 960.085 4.255 960.415 4.270 ;
        RECT 995.965 4.255 996.295 4.270 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.850 14.010 1012.990 15.300 ;
        RECT 1012.620 13.870 1012.990 14.010 ;
        RECT 1012.620 6.645 1012.760 13.870 ;
        RECT 978.050 6.275 978.330 6.645 ;
        RECT 1012.550 6.275 1012.830 6.645 ;
        RECT 978.120 2.400 978.260 6.275 ;
        RECT 977.910 -4.800 978.470 2.400 ;
      LAYER met3 ;
        RECT 978.025 6.610 978.355 6.625 ;
        RECT 1012.525 6.610 1012.855 6.625 ;
        RECT 978.025 6.310 1012.855 6.610 ;
        RECT 978.025 6.295 978.355 6.310 ;
        RECT 1012.525 6.295 1012.855 6.310 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 660.170 6.700 660.490 6.760 ;
        RECT 714.450 6.700 714.770 6.760 ;
        RECT 660.170 6.560 714.770 6.700 ;
        RECT 660.170 6.500 660.490 6.560 ;
        RECT 714.450 6.500 714.770 6.560 ;
      LAYER met2 ;
        RECT 714.770 14.010 714.910 15.300 ;
        RECT 714.540 13.870 714.910 14.010 ;
        RECT 714.540 6.790 714.680 13.870 ;
        RECT 660.200 6.470 660.460 6.790 ;
        RECT 714.480 6.470 714.740 6.790 ;
        RECT 660.260 3.810 660.400 6.470 ;
        RECT 658.880 3.670 660.400 3.810 ;
        RECT 658.880 2.400 659.020 3.670 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.410 14.010 1029.550 15.300 ;
        RECT 1029.180 13.870 1029.550 14.010 ;
        RECT 1029.180 3.925 1029.320 13.870 ;
        RECT 995.530 3.555 995.810 3.925 ;
        RECT 1029.110 3.555 1029.390 3.925 ;
        RECT 995.600 2.400 995.740 3.555 ;
        RECT 995.390 -4.800 995.950 2.400 ;
      LAYER met3 ;
        RECT 995.505 3.890 995.835 3.905 ;
        RECT 1029.085 3.890 1029.415 3.905 ;
        RECT 995.505 3.590 1029.415 3.890 ;
        RECT 995.505 3.575 995.835 3.590 ;
        RECT 1029.085 3.575 1029.415 3.590 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.970 14.010 1046.110 15.300 ;
        RECT 1045.740 13.870 1046.110 14.010 ;
        RECT 1045.740 5.285 1045.880 13.870 ;
        RECT 1013.470 4.915 1013.750 5.285 ;
        RECT 1045.670 4.915 1045.950 5.285 ;
        RECT 1013.540 2.400 1013.680 4.915 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER met3 ;
        RECT 1013.445 5.250 1013.775 5.265 ;
        RECT 1045.645 5.250 1045.975 5.265 ;
        RECT 1013.445 4.950 1045.975 5.250 ;
        RECT 1013.445 4.935 1013.775 4.950 ;
        RECT 1045.645 4.935 1045.975 4.950 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.530 14.010 1062.670 15.300 ;
        RECT 1062.300 13.870 1062.670 14.010 ;
        RECT 1062.300 8.005 1062.440 13.870 ;
        RECT 1030.950 7.635 1031.230 8.005 ;
        RECT 1062.230 7.635 1062.510 8.005 ;
        RECT 1031.020 2.400 1031.160 7.635 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
      LAYER met3 ;
        RECT 1030.925 7.970 1031.255 7.985 ;
        RECT 1062.205 7.970 1062.535 7.985 ;
        RECT 1030.925 7.670 1062.535 7.970 ;
        RECT 1030.925 7.655 1031.255 7.670 ;
        RECT 1062.205 7.655 1062.535 7.670 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.090 14.010 1079.230 15.300 ;
        RECT 1078.860 13.870 1079.230 14.010 ;
        RECT 1078.860 11.405 1079.000 13.870 ;
        RECT 1048.890 11.035 1049.170 11.405 ;
        RECT 1078.790 11.035 1079.070 11.405 ;
        RECT 1048.960 2.400 1049.100 11.035 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
      LAYER met3 ;
        RECT 1048.865 11.370 1049.195 11.385 ;
        RECT 1078.765 11.370 1079.095 11.385 ;
        RECT 1048.865 11.070 1079.095 11.370 ;
        RECT 1048.865 11.055 1049.195 11.070 ;
        RECT 1078.765 11.055 1079.095 11.070 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.650 14.010 1095.790 15.300 ;
        RECT 1095.420 13.870 1095.790 14.010 ;
        RECT 1095.420 8.685 1095.560 13.870 ;
        RECT 1066.830 8.315 1067.110 8.685 ;
        RECT 1095.350 8.315 1095.630 8.685 ;
        RECT 1066.900 2.400 1067.040 8.315 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
      LAYER met3 ;
        RECT 1066.805 8.650 1067.135 8.665 ;
        RECT 1095.325 8.650 1095.655 8.665 ;
        RECT 1066.805 8.350 1095.655 8.650 ;
        RECT 1066.805 8.335 1067.135 8.350 ;
        RECT 1095.325 8.335 1095.655 8.350 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.210 14.010 1112.350 15.300 ;
        RECT 1111.980 13.870 1112.350 14.010 ;
        RECT 1111.980 12.085 1112.120 13.870 ;
        RECT 1084.310 11.715 1084.590 12.085 ;
        RECT 1111.910 11.715 1112.190 12.085 ;
        RECT 1084.380 2.400 1084.520 11.715 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
      LAYER met3 ;
        RECT 1084.285 12.050 1084.615 12.065 ;
        RECT 1111.885 12.050 1112.215 12.065 ;
        RECT 1084.285 11.750 1112.215 12.050 ;
        RECT 1084.285 11.735 1084.615 11.750 ;
        RECT 1111.885 11.735 1112.215 11.750 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.770 14.010 1128.910 15.300 ;
        RECT 1128.540 13.870 1128.910 14.010 ;
        RECT 1128.540 10.045 1128.680 13.870 ;
        RECT 1102.250 9.675 1102.530 10.045 ;
        RECT 1128.470 9.675 1128.750 10.045 ;
        RECT 1102.320 2.400 1102.460 9.675 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
      LAYER met3 ;
        RECT 1102.225 10.010 1102.555 10.025 ;
        RECT 1128.445 10.010 1128.775 10.025 ;
        RECT 1102.225 9.710 1128.775 10.010 ;
        RECT 1102.225 9.695 1102.555 9.710 ;
        RECT 1128.445 9.695 1128.775 9.710 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.330 14.010 1145.470 15.300 ;
        RECT 1145.100 13.870 1145.470 14.010 ;
        RECT 1145.100 10.725 1145.240 13.870 ;
        RECT 1119.730 10.355 1120.010 10.725 ;
        RECT 1145.030 10.355 1145.310 10.725 ;
        RECT 1119.800 2.400 1119.940 10.355 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
      LAYER met3 ;
        RECT 1119.705 10.690 1120.035 10.705 ;
        RECT 1145.005 10.690 1145.335 10.705 ;
        RECT 1119.705 10.390 1145.335 10.690 ;
        RECT 1119.705 10.375 1120.035 10.390 ;
        RECT 1145.005 10.375 1145.335 10.390 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.890 14.010 1162.030 15.300 ;
        RECT 1161.660 13.870 1162.030 14.010 ;
        RECT 1161.660 10.045 1161.800 13.870 ;
        RECT 1137.670 9.675 1137.950 10.045 ;
        RECT 1161.590 9.675 1161.870 10.045 ;
        RECT 1137.740 2.400 1137.880 9.675 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
      LAYER met3 ;
        RECT 1137.645 10.010 1137.975 10.025 ;
        RECT 1161.565 10.010 1161.895 10.025 ;
        RECT 1137.645 9.710 1161.895 10.010 ;
        RECT 1137.645 9.695 1137.975 9.710 ;
        RECT 1161.565 9.695 1161.895 9.710 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.450 14.010 1178.590 15.300 ;
        RECT 1178.220 13.870 1178.590 14.010 ;
        RECT 1178.220 7.325 1178.360 13.870 ;
        RECT 1155.150 6.955 1155.430 7.325 ;
        RECT 1178.150 6.955 1178.430 7.325 ;
        RECT 1155.220 2.400 1155.360 6.955 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
      LAYER met3 ;
        RECT 1155.125 7.290 1155.455 7.305 ;
        RECT 1178.125 7.290 1178.455 7.305 ;
        RECT 1155.125 6.990 1178.455 7.290 ;
        RECT 1155.125 6.975 1155.455 6.990 ;
        RECT 1178.125 6.975 1178.455 6.990 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.330 14.010 731.470 15.300 ;
        RECT 731.100 13.870 731.470 14.010 ;
        RECT 731.100 10.045 731.240 13.870 ;
        RECT 676.290 9.675 676.570 10.045 ;
        RECT 731.030 9.675 731.310 10.045 ;
        RECT 676.360 2.400 676.500 9.675 ;
        RECT 676.150 -4.800 676.710 2.400 ;
      LAYER met3 ;
        RECT 676.265 10.010 676.595 10.025 ;
        RECT 731.005 10.010 731.335 10.025 ;
        RECT 676.265 9.710 731.335 10.010 ;
        RECT 676.265 9.695 676.595 9.710 ;
        RECT 731.005 9.695 731.335 9.710 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.010 14.010 1195.150 15.300 ;
        RECT 1194.780 13.870 1195.150 14.010 ;
        RECT 1194.780 8.685 1194.920 13.870 ;
        RECT 1173.090 8.315 1173.370 8.685 ;
        RECT 1194.710 8.315 1194.990 8.685 ;
        RECT 1173.160 2.400 1173.300 8.315 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
      LAYER met3 ;
        RECT 1173.065 8.650 1173.395 8.665 ;
        RECT 1194.685 8.650 1195.015 8.665 ;
        RECT 1173.065 8.350 1195.015 8.650 ;
        RECT 1173.065 8.335 1173.395 8.350 ;
        RECT 1194.685 8.335 1195.015 8.350 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.570 14.010 1211.710 15.300 ;
        RECT 1211.340 13.870 1211.710 14.010 ;
        RECT 1211.340 10.045 1211.480 13.870 ;
        RECT 1190.570 9.675 1190.850 10.045 ;
        RECT 1211.270 9.675 1211.550 10.045 ;
        RECT 1190.640 2.400 1190.780 9.675 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
      LAYER met3 ;
        RECT 1190.545 10.010 1190.875 10.025 ;
        RECT 1211.245 10.010 1211.575 10.025 ;
        RECT 1190.545 9.710 1211.575 10.010 ;
        RECT 1190.545 9.695 1190.875 9.710 ;
        RECT 1211.245 9.695 1211.575 9.710 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.130 14.010 1228.270 15.300 ;
        RECT 1227.900 13.870 1228.270 14.010 ;
        RECT 1227.900 9.365 1228.040 13.870 ;
        RECT 1208.510 8.995 1208.790 9.365 ;
        RECT 1227.830 8.995 1228.110 9.365 ;
        RECT 1208.580 2.400 1208.720 8.995 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
      LAYER met3 ;
        RECT 1208.485 9.330 1208.815 9.345 ;
        RECT 1227.805 9.330 1228.135 9.345 ;
        RECT 1208.485 9.030 1228.135 9.330 ;
        RECT 1208.485 9.015 1208.815 9.030 ;
        RECT 1227.805 9.015 1228.135 9.030 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.690 14.010 1244.830 15.300 ;
        RECT 1244.460 13.870 1244.830 14.010 ;
        RECT 1244.460 7.325 1244.600 13.870 ;
        RECT 1225.990 6.955 1226.270 7.325 ;
        RECT 1244.390 6.955 1244.670 7.325 ;
        RECT 1226.060 2.400 1226.200 6.955 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
      LAYER met3 ;
        RECT 1225.965 7.290 1226.295 7.305 ;
        RECT 1244.365 7.290 1244.695 7.305 ;
        RECT 1225.965 6.990 1244.695 7.290 ;
        RECT 1225.965 6.975 1226.295 6.990 ;
        RECT 1244.365 6.975 1244.695 6.990 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.250 14.010 1261.390 15.300 ;
        RECT 1261.020 13.870 1261.390 14.010 ;
        RECT 1261.020 10.045 1261.160 13.870 ;
        RECT 1243.930 9.675 1244.210 10.045 ;
        RECT 1260.950 9.675 1261.230 10.045 ;
        RECT 1244.000 2.400 1244.140 9.675 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
      LAYER met3 ;
        RECT 1243.905 10.010 1244.235 10.025 ;
        RECT 1260.925 10.010 1261.255 10.025 ;
        RECT 1243.905 9.710 1261.255 10.010 ;
        RECT 1243.905 9.695 1244.235 9.710 ;
        RECT 1260.925 9.695 1261.255 9.710 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.810 14.010 1277.950 15.300 ;
        RECT 1277.580 13.870 1277.950 14.010 ;
        RECT 1277.580 7.325 1277.720 13.870 ;
        RECT 1261.870 6.955 1262.150 7.325 ;
        RECT 1277.510 6.955 1277.790 7.325 ;
        RECT 1261.940 2.400 1262.080 6.955 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
      LAYER met3 ;
        RECT 1261.845 7.290 1262.175 7.305 ;
        RECT 1277.485 7.290 1277.815 7.305 ;
        RECT 1261.845 6.990 1277.815 7.290 ;
        RECT 1261.845 6.975 1262.175 6.990 ;
        RECT 1277.485 6.975 1277.815 6.990 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.370 14.010 1294.510 15.300 ;
        RECT 1294.140 13.870 1294.510 14.010 ;
        RECT 1294.140 7.325 1294.280 13.870 ;
        RECT 1279.350 6.955 1279.630 7.325 ;
        RECT 1294.070 6.955 1294.350 7.325 ;
        RECT 1279.420 2.400 1279.560 6.955 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
      LAYER met3 ;
        RECT 1279.325 7.290 1279.655 7.305 ;
        RECT 1294.045 7.290 1294.375 7.305 ;
        RECT 1279.325 6.990 1294.375 7.290 ;
        RECT 1279.325 6.975 1279.655 6.990 ;
        RECT 1294.045 6.975 1294.375 6.990 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.930 14.010 1311.070 15.300 ;
        RECT 1310.700 13.870 1311.070 14.010 ;
        RECT 1310.700 6.645 1310.840 13.870 ;
        RECT 1297.290 6.275 1297.570 6.645 ;
        RECT 1310.630 6.275 1310.910 6.645 ;
        RECT 1297.360 2.400 1297.500 6.275 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
      LAYER met3 ;
        RECT 1297.265 6.610 1297.595 6.625 ;
        RECT 1310.605 6.610 1310.935 6.625 ;
        RECT 1297.265 6.310 1310.935 6.610 ;
        RECT 1297.265 6.295 1297.595 6.310 ;
        RECT 1310.605 6.295 1310.935 6.310 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.490 14.010 1327.630 15.300 ;
        RECT 1327.260 13.870 1327.630 14.010 ;
        RECT 1327.260 7.325 1327.400 13.870 ;
        RECT 1314.770 6.955 1315.050 7.325 ;
        RECT 1327.190 6.955 1327.470 7.325 ;
        RECT 1314.840 2.400 1314.980 6.955 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
      LAYER met3 ;
        RECT 1314.745 7.290 1315.075 7.305 ;
        RECT 1327.165 7.290 1327.495 7.305 ;
        RECT 1314.745 6.990 1327.495 7.290 ;
        RECT 1314.745 6.975 1315.075 6.990 ;
        RECT 1327.165 6.975 1327.495 6.990 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.050 14.010 1344.190 15.300 ;
        RECT 1343.820 13.870 1344.190 14.010 ;
        RECT 1343.820 5.965 1343.960 13.870 ;
        RECT 1332.710 5.595 1332.990 5.965 ;
        RECT 1343.750 5.595 1344.030 5.965 ;
        RECT 1332.780 2.400 1332.920 5.595 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
      LAYER met3 ;
        RECT 1332.685 5.930 1333.015 5.945 ;
        RECT 1343.725 5.930 1344.055 5.945 ;
        RECT 1332.685 5.630 1344.055 5.930 ;
        RECT 1332.685 5.615 1333.015 5.630 ;
        RECT 1343.725 5.615 1344.055 5.630 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.050 0.580 696.370 0.640 ;
        RECT 746.650 0.580 746.970 0.640 ;
        RECT 696.050 0.440 746.970 0.580 ;
        RECT 696.050 0.380 696.370 0.440 ;
        RECT 746.650 0.380 746.970 0.440 ;
      LAYER met2 ;
        RECT 747.890 14.010 748.030 15.300 ;
        RECT 746.740 13.870 748.030 14.010 ;
        RECT 694.090 0.410 694.650 2.400 ;
        RECT 746.740 0.670 746.880 13.870 ;
        RECT 696.080 0.410 696.340 0.670 ;
        RECT 694.090 0.350 696.340 0.410 ;
        RECT 746.680 0.350 746.940 0.670 ;
        RECT 694.090 0.270 696.280 0.350 ;
        RECT 694.090 -4.800 694.650 0.270 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.610 14.010 1360.750 15.300 ;
        RECT 1360.380 13.870 1360.750 14.010 ;
        RECT 1360.380 8.005 1360.520 13.870 ;
        RECT 1350.190 7.635 1350.470 8.005 ;
        RECT 1360.310 7.635 1360.590 8.005 ;
        RECT 1350.260 2.400 1350.400 7.635 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
      LAYER met3 ;
        RECT 1350.165 7.970 1350.495 7.985 ;
        RECT 1360.285 7.970 1360.615 7.985 ;
        RECT 1350.165 7.670 1360.615 7.970 ;
        RECT 1350.165 7.655 1350.495 7.670 ;
        RECT 1360.285 7.655 1360.615 7.670 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.170 14.010 1377.310 15.300 ;
        RECT 1376.940 13.870 1377.310 14.010 ;
        RECT 1376.940 6.645 1377.080 13.870 ;
        RECT 1368.130 6.275 1368.410 6.645 ;
        RECT 1376.870 6.275 1377.150 6.645 ;
        RECT 1368.200 2.400 1368.340 6.275 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
      LAYER met3 ;
        RECT 1368.105 6.610 1368.435 6.625 ;
        RECT 1376.845 6.610 1377.175 6.625 ;
        RECT 1368.105 6.310 1377.175 6.610 ;
        RECT 1368.105 6.295 1368.435 6.310 ;
        RECT 1376.845 6.295 1377.175 6.310 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.730 14.010 1393.870 15.300 ;
        RECT 1393.500 13.870 1393.870 14.010 ;
        RECT 1393.500 5.965 1393.640 13.870 ;
        RECT 1385.610 5.595 1385.890 5.965 ;
        RECT 1393.430 5.595 1393.710 5.965 ;
        RECT 1385.680 2.400 1385.820 5.595 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
      LAYER met3 ;
        RECT 1385.585 5.930 1385.915 5.945 ;
        RECT 1393.405 5.930 1393.735 5.945 ;
        RECT 1385.585 5.630 1393.735 5.930 ;
        RECT 1385.585 5.615 1385.915 5.630 ;
        RECT 1393.405 5.615 1393.735 5.630 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.290 14.010 1410.430 15.300 ;
        RECT 1410.060 13.870 1410.430 14.010 ;
        RECT 1410.060 5.965 1410.200 13.870 ;
        RECT 1403.550 5.595 1403.830 5.965 ;
        RECT 1409.990 5.595 1410.270 5.965 ;
        RECT 1403.620 2.400 1403.760 5.595 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
      LAYER met3 ;
        RECT 1403.525 5.930 1403.855 5.945 ;
        RECT 1409.965 5.930 1410.295 5.945 ;
        RECT 1403.525 5.630 1410.295 5.930 ;
        RECT 1403.525 5.615 1403.855 5.630 ;
        RECT 1409.965 5.615 1410.295 5.630 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.850 14.010 1426.990 15.300 ;
        RECT 1421.560 13.870 1426.990 14.010 ;
        RECT 1421.560 2.400 1421.700 13.870 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.410 14.010 1443.550 15.300 ;
        RECT 1443.180 13.870 1443.550 14.010 ;
        RECT 1443.180 6.645 1443.320 13.870 ;
        RECT 1438.970 6.275 1439.250 6.645 ;
        RECT 1443.110 6.275 1443.390 6.645 ;
        RECT 1439.040 2.400 1439.180 6.275 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
      LAYER met3 ;
        RECT 1438.945 6.610 1439.275 6.625 ;
        RECT 1443.085 6.610 1443.415 6.625 ;
        RECT 1438.945 6.310 1443.415 6.610 ;
        RECT 1438.945 6.295 1439.275 6.310 ;
        RECT 1443.085 6.295 1443.415 6.310 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.970 14.010 1460.110 15.300 ;
        RECT 1459.280 13.870 1460.110 14.010 ;
        RECT 1456.770 1.770 1457.330 2.400 ;
        RECT 1459.280 1.770 1459.420 13.870 ;
        RECT 1456.770 1.630 1459.420 1.770 ;
        RECT 1456.770 -4.800 1457.330 1.630 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.530 14.010 1476.670 15.300 ;
        RECT 1476.300 13.870 1476.670 14.010 ;
        RECT 1474.250 1.770 1474.810 2.400 ;
        RECT 1476.300 1.770 1476.440 13.870 ;
        RECT 1474.250 1.630 1476.440 1.770 ;
        RECT 1474.250 -4.800 1474.810 1.630 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.090 14.010 1493.230 15.300 ;
        RECT 1492.400 13.870 1493.230 14.010 ;
        RECT 1492.400 2.400 1492.540 13.870 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.650 14.010 1509.790 15.300 ;
        RECT 1509.650 13.870 1510.020 14.010 ;
        RECT 1509.880 2.400 1510.020 13.870 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.450 14.010 764.590 15.300 ;
        RECT 764.220 13.870 764.590 14.010 ;
        RECT 764.220 10.725 764.360 13.870 ;
        RECT 712.170 10.355 712.450 10.725 ;
        RECT 764.150 10.355 764.430 10.725 ;
        RECT 712.240 2.400 712.380 10.355 ;
        RECT 712.030 -4.800 712.590 2.400 ;
      LAYER met3 ;
        RECT 712.145 10.690 712.475 10.705 ;
        RECT 764.125 10.690 764.455 10.705 ;
        RECT 712.145 10.390 764.455 10.690 ;
        RECT 712.145 10.375 712.475 10.390 ;
        RECT 764.125 10.375 764.455 10.390 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.210 14.010 1526.350 15.300 ;
        RECT 1526.210 13.870 1527.960 14.010 ;
        RECT 1527.820 2.400 1527.960 13.870 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.770 14.010 1542.910 15.300 ;
        RECT 1542.770 13.870 1545.440 14.010 ;
        RECT 1545.300 2.400 1545.440 13.870 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.330 14.010 1559.470 15.300 ;
        RECT 1559.330 13.870 1561.080 14.010 ;
        RECT 1560.940 1.770 1561.080 13.870 ;
        RECT 1563.030 1.770 1563.590 2.400 ;
        RECT 1560.940 1.630 1563.590 1.770 ;
        RECT 1563.030 -4.800 1563.590 1.630 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.890 14.010 1576.030 15.300 ;
        RECT 1575.890 13.870 1576.260 14.010 ;
        RECT 1576.120 6.645 1576.260 13.870 ;
        RECT 1576.050 6.275 1576.330 6.645 ;
        RECT 1581.110 6.275 1581.390 6.645 ;
        RECT 1581.180 2.400 1581.320 6.275 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
      LAYER met3 ;
        RECT 1576.025 6.610 1576.355 6.625 ;
        RECT 1581.085 6.610 1581.415 6.625 ;
        RECT 1576.025 6.310 1581.415 6.610 ;
        RECT 1576.025 6.295 1576.355 6.310 ;
        RECT 1581.085 6.295 1581.415 6.310 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.450 14.010 1592.590 15.300 ;
        RECT 1592.220 13.870 1592.590 14.010 ;
        RECT 1592.220 5.965 1592.360 13.870 ;
        RECT 1592.150 5.595 1592.430 5.965 ;
        RECT 1598.590 5.595 1598.870 5.965 ;
        RECT 1598.660 2.400 1598.800 5.595 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
      LAYER met3 ;
        RECT 1592.125 5.930 1592.455 5.945 ;
        RECT 1598.565 5.930 1598.895 5.945 ;
        RECT 1592.125 5.630 1598.895 5.930 ;
        RECT 1592.125 5.615 1592.455 5.630 ;
        RECT 1598.565 5.615 1598.895 5.630 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.010 14.010 1609.150 15.300 ;
        RECT 1609.010 13.870 1609.380 14.010 ;
        RECT 1609.240 5.285 1609.380 13.870 ;
        RECT 1609.170 4.915 1609.450 5.285 ;
        RECT 1616.530 4.915 1616.810 5.285 ;
        RECT 1616.600 2.400 1616.740 4.915 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
      LAYER met3 ;
        RECT 1609.145 5.250 1609.475 5.265 ;
        RECT 1616.505 5.250 1616.835 5.265 ;
        RECT 1609.145 4.950 1616.835 5.250 ;
        RECT 1609.145 4.935 1609.475 4.950 ;
        RECT 1616.505 4.935 1616.835 4.950 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.570 14.010 1625.710 15.300 ;
        RECT 1625.570 13.870 1625.940 14.010 ;
        RECT 1625.800 6.645 1625.940 13.870 ;
        RECT 1625.730 6.275 1626.010 6.645 ;
        RECT 1634.010 6.275 1634.290 6.645 ;
        RECT 1634.080 2.400 1634.220 6.275 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
      LAYER met3 ;
        RECT 1625.705 6.610 1626.035 6.625 ;
        RECT 1633.985 6.610 1634.315 6.625 ;
        RECT 1625.705 6.310 1634.315 6.610 ;
        RECT 1625.705 6.295 1626.035 6.310 ;
        RECT 1633.985 6.295 1634.315 6.310 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.130 14.010 1642.270 15.300 ;
        RECT 1641.900 13.870 1642.270 14.010 ;
        RECT 1641.900 5.965 1642.040 13.870 ;
        RECT 1641.830 5.595 1642.110 5.965 ;
        RECT 1651.950 5.595 1652.230 5.965 ;
        RECT 1652.020 2.400 1652.160 5.595 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
      LAYER met3 ;
        RECT 1641.805 5.930 1642.135 5.945 ;
        RECT 1651.925 5.930 1652.255 5.945 ;
        RECT 1641.805 5.630 1652.255 5.930 ;
        RECT 1641.805 5.615 1642.135 5.630 ;
        RECT 1651.925 5.615 1652.255 5.630 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.690 14.010 1658.830 15.300 ;
        RECT 1658.690 13.870 1659.060 14.010 ;
        RECT 1658.920 4.605 1659.060 13.870 ;
        RECT 1658.850 4.235 1659.130 4.605 ;
        RECT 1669.430 4.235 1669.710 4.605 ;
        RECT 1669.500 2.400 1669.640 4.235 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
      LAYER met3 ;
        RECT 1658.825 4.570 1659.155 4.585 ;
        RECT 1669.405 4.570 1669.735 4.585 ;
        RECT 1658.825 4.270 1669.735 4.570 ;
        RECT 1658.825 4.255 1659.155 4.270 ;
        RECT 1669.405 4.255 1669.735 4.270 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.250 14.010 1675.390 15.300 ;
        RECT 1675.250 13.870 1675.620 14.010 ;
        RECT 1675.480 6.645 1675.620 13.870 ;
        RECT 1675.410 6.275 1675.690 6.645 ;
        RECT 1687.370 6.275 1687.650 6.645 ;
        RECT 1687.440 2.400 1687.580 6.275 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
      LAYER met3 ;
        RECT 1675.385 6.610 1675.715 6.625 ;
        RECT 1687.345 6.610 1687.675 6.625 ;
        RECT 1675.385 6.310 1687.675 6.610 ;
        RECT 1675.385 6.295 1675.715 6.310 ;
        RECT 1687.345 6.295 1687.675 6.310 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.010 6.700 731.330 6.760 ;
        RECT 780.690 6.700 781.010 6.760 ;
        RECT 731.010 6.560 781.010 6.700 ;
        RECT 731.010 6.500 731.330 6.560 ;
        RECT 780.690 6.500 781.010 6.560 ;
      LAYER met2 ;
        RECT 781.010 14.010 781.150 15.300 ;
        RECT 780.780 13.870 781.150 14.010 ;
        RECT 780.780 6.790 780.920 13.870 ;
        RECT 731.040 6.470 731.300 6.790 ;
        RECT 780.720 6.470 780.980 6.790 ;
        RECT 731.100 3.810 731.240 6.470 ;
        RECT 729.720 3.670 731.240 3.810 ;
        RECT 729.720 2.400 729.860 3.670 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.810 14.010 1691.950 15.300 ;
        RECT 1691.810 13.870 1692.180 14.010 ;
        RECT 1692.040 6.645 1692.180 13.870 ;
        RECT 1691.970 6.275 1692.250 6.645 ;
        RECT 1704.850 6.275 1705.130 6.645 ;
        RECT 1704.920 2.400 1705.060 6.275 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
      LAYER met3 ;
        RECT 1691.945 6.610 1692.275 6.625 ;
        RECT 1704.825 6.610 1705.155 6.625 ;
        RECT 1691.945 6.310 1705.155 6.610 ;
        RECT 1691.945 6.295 1692.275 6.310 ;
        RECT 1704.825 6.295 1705.155 6.310 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.370 14.010 1708.510 15.300 ;
        RECT 1708.370 13.870 1708.740 14.010 ;
        RECT 1708.600 6.645 1708.740 13.870 ;
        RECT 1708.530 6.275 1708.810 6.645 ;
        RECT 1722.790 6.275 1723.070 6.645 ;
        RECT 1722.860 2.400 1723.000 6.275 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
      LAYER met3 ;
        RECT 1708.505 6.610 1708.835 6.625 ;
        RECT 1722.765 6.610 1723.095 6.625 ;
        RECT 1708.505 6.310 1723.095 6.610 ;
        RECT 1708.505 6.295 1708.835 6.310 ;
        RECT 1722.765 6.295 1723.095 6.310 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.930 14.125 1725.070 15.300 ;
        RECT 1724.860 13.755 1725.140 14.125 ;
        RECT 1738.890 13.330 1739.170 13.445 ;
        RECT 1738.890 13.190 1740.480 13.330 ;
        RECT 1738.890 13.075 1739.170 13.190 ;
        RECT 1740.340 2.400 1740.480 13.190 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
      LAYER met3 ;
        RECT 1724.835 14.090 1725.165 14.105 ;
        RECT 1724.835 13.790 1729.290 14.090 ;
        RECT 1724.835 13.775 1725.165 13.790 ;
        RECT 1728.990 13.410 1729.290 13.790 ;
        RECT 1738.865 13.410 1739.195 13.425 ;
        RECT 1728.990 13.110 1739.195 13.410 ;
        RECT 1738.865 13.095 1739.195 13.110 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.490 14.010 1741.630 15.300 ;
        RECT 1741.490 13.870 1741.860 14.010 ;
        RECT 1741.720 5.965 1741.860 13.870 ;
        RECT 1741.650 5.595 1741.930 5.965 ;
        RECT 1758.210 5.595 1758.490 5.965 ;
        RECT 1758.280 2.400 1758.420 5.595 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
      LAYER met3 ;
        RECT 1741.625 5.930 1741.955 5.945 ;
        RECT 1758.185 5.930 1758.515 5.945 ;
        RECT 1741.625 5.630 1758.515 5.930 ;
        RECT 1741.625 5.615 1741.955 5.630 ;
        RECT 1758.185 5.615 1758.515 5.630 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1757.960 14.180 1758.280 14.240 ;
        RECT 1775.210 14.180 1775.530 14.240 ;
        RECT 1757.960 14.040 1775.530 14.180 ;
        RECT 1757.960 13.980 1758.280 14.040 ;
        RECT 1775.210 13.980 1775.530 14.040 ;
      LAYER met2 ;
        RECT 1758.050 14.270 1758.190 15.300 ;
        RECT 1757.990 13.950 1758.250 14.270 ;
        RECT 1775.240 13.950 1775.500 14.270 ;
        RECT 1775.300 7.210 1775.440 13.950 ;
        RECT 1775.300 7.070 1776.360 7.210 ;
        RECT 1776.220 2.400 1776.360 7.070 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.610 14.010 1774.750 15.300 ;
        RECT 1774.610 13.870 1774.980 14.010 ;
        RECT 1774.840 6.645 1774.980 13.870 ;
        RECT 1774.770 6.275 1775.050 6.645 ;
        RECT 1793.630 6.275 1793.910 6.645 ;
        RECT 1793.700 2.400 1793.840 6.275 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
      LAYER met3 ;
        RECT 1774.745 6.610 1775.075 6.625 ;
        RECT 1793.605 6.610 1793.935 6.625 ;
        RECT 1774.745 6.310 1793.935 6.610 ;
        RECT 1774.745 6.295 1775.075 6.310 ;
        RECT 1793.605 6.295 1793.935 6.310 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1791.080 14.180 1791.400 14.240 ;
        RECT 1808.330 14.180 1808.650 14.240 ;
        RECT 1791.080 14.040 1808.650 14.180 ;
        RECT 1791.080 13.980 1791.400 14.040 ;
        RECT 1808.330 13.980 1808.650 14.040 ;
      LAYER met2 ;
        RECT 1791.170 14.270 1791.310 15.300 ;
        RECT 1791.110 13.950 1791.370 14.270 ;
        RECT 1808.360 14.010 1808.620 14.270 ;
        RECT 1808.360 13.950 1809.480 14.010 ;
        RECT 1808.420 13.870 1809.480 13.950 ;
        RECT 1809.340 1.770 1809.480 13.870 ;
        RECT 1811.430 1.770 1811.990 2.400 ;
        RECT 1809.340 1.630 1811.990 1.770 ;
        RECT 1811.430 -4.800 1811.990 1.630 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1820.290 14.520 1820.610 14.580 ;
        RECT 1828.570 14.520 1828.890 14.580 ;
        RECT 1820.290 14.380 1828.890 14.520 ;
        RECT 1820.290 14.320 1820.610 14.380 ;
        RECT 1828.570 14.320 1828.890 14.380 ;
      LAYER met2 ;
        RECT 1807.730 14.125 1807.870 15.300 ;
        RECT 1820.320 14.290 1820.580 14.610 ;
        RECT 1828.600 14.290 1828.860 14.610 ;
        RECT 1820.380 14.125 1820.520 14.290 ;
        RECT 1807.660 13.755 1807.940 14.125 ;
        RECT 1820.310 13.755 1820.590 14.125 ;
        RECT 1828.660 7.210 1828.800 14.290 ;
        RECT 1828.660 7.070 1829.260 7.210 ;
        RECT 1829.120 2.400 1829.260 7.070 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
      LAYER met3 ;
        RECT 1807.635 14.090 1807.965 14.105 ;
        RECT 1820.285 14.090 1820.615 14.105 ;
        RECT 1807.635 13.790 1820.615 14.090 ;
        RECT 1807.635 13.775 1807.965 13.790 ;
        RECT 1820.285 13.775 1820.615 13.790 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.290 14.125 1824.430 15.300 ;
        RECT 1824.220 13.755 1824.500 14.125 ;
        RECT 1845.150 13.330 1845.430 13.445 ;
        RECT 1845.150 13.190 1847.200 13.330 ;
        RECT 1845.150 13.075 1845.430 13.190 ;
        RECT 1847.060 2.400 1847.200 13.190 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
      LAYER met3 ;
        RECT 1824.195 14.090 1824.525 14.105 ;
        RECT 1824.195 13.790 1839.690 14.090 ;
        RECT 1824.195 13.775 1824.525 13.790 ;
        RECT 1839.390 13.410 1839.690 13.790 ;
        RECT 1845.125 13.410 1845.455 13.425 ;
        RECT 1839.390 13.110 1845.455 13.410 ;
        RECT 1845.125 13.095 1845.455 13.110 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1841.450 7.720 1841.770 7.780 ;
        RECT 1863.070 7.720 1863.390 7.780 ;
        RECT 1841.450 7.580 1863.390 7.720 ;
        RECT 1841.450 7.520 1841.770 7.580 ;
        RECT 1863.070 7.520 1863.390 7.580 ;
      LAYER met2 ;
        RECT 1840.850 14.690 1840.990 15.300 ;
        RECT 1840.850 14.550 1841.680 14.690 ;
        RECT 1841.540 7.810 1841.680 14.550 ;
        RECT 1841.480 7.490 1841.740 7.810 ;
        RECT 1863.100 7.490 1863.360 7.810 ;
        RECT 1863.160 7.210 1863.300 7.490 ;
        RECT 1863.160 7.070 1864.680 7.210 ;
        RECT 1864.540 2.400 1864.680 7.070 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.570 14.010 797.710 15.300 ;
        RECT 797.340 13.870 797.710 14.010 ;
        RECT 797.340 12.765 797.480 13.870 ;
        RECT 747.590 12.395 747.870 12.765 ;
        RECT 797.270 12.395 797.550 12.765 ;
        RECT 747.660 2.400 747.800 12.395 ;
        RECT 747.450 -4.800 748.010 2.400 ;
      LAYER met3 ;
        RECT 747.565 12.730 747.895 12.745 ;
        RECT 797.245 12.730 797.575 12.745 ;
        RECT 747.565 12.430 797.575 12.730 ;
        RECT 747.565 12.415 747.895 12.430 ;
        RECT 797.245 12.415 797.575 12.430 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.410 14.125 1857.550 15.300 ;
        RECT 1857.340 13.755 1857.620 14.125 ;
        RECT 1882.410 13.755 1882.690 14.125 ;
        RECT 1882.480 2.400 1882.620 13.755 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
      LAYER met3 ;
        RECT 1857.315 14.090 1857.645 14.105 ;
        RECT 1882.385 14.090 1882.715 14.105 ;
        RECT 1857.315 13.790 1861.770 14.090 ;
        RECT 1857.315 13.775 1857.645 13.790 ;
        RECT 1861.470 13.410 1861.770 13.790 ;
        RECT 1864.230 13.790 1882.715 14.090 ;
        RECT 1864.230 13.410 1864.530 13.790 ;
        RECT 1882.385 13.775 1882.715 13.790 ;
        RECT 1861.470 13.110 1864.530 13.410 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.970 14.010 1874.110 15.300 ;
        RECT 1873.970 13.870 1874.340 14.010 ;
        RECT 1874.200 13.445 1874.340 13.870 ;
        RECT 1874.130 13.075 1874.410 13.445 ;
        RECT 1897.590 13.075 1897.870 13.445 ;
        RECT 1897.660 1.770 1897.800 13.075 ;
        RECT 1899.750 1.770 1900.310 2.400 ;
        RECT 1897.660 1.630 1900.310 1.770 ;
        RECT 1899.750 -4.800 1900.310 1.630 ;
      LAYER met3 ;
        RECT 1883.550 13.790 1893.050 14.090 ;
        RECT 1874.105 13.410 1874.435 13.425 ;
        RECT 1883.550 13.410 1883.850 13.790 ;
        RECT 1874.105 13.110 1883.850 13.410 ;
        RECT 1892.750 13.410 1893.050 13.790 ;
        RECT 1897.565 13.410 1897.895 13.425 ;
        RECT 1892.750 13.110 1897.895 13.410 ;
        RECT 1874.105 13.095 1874.435 13.110 ;
        RECT 1897.565 13.095 1897.895 13.110 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1890.670 13.840 1890.990 13.900 ;
        RECT 1917.350 13.840 1917.670 13.900 ;
        RECT 1890.670 13.700 1917.670 13.840 ;
        RECT 1890.670 13.640 1890.990 13.700 ;
        RECT 1917.350 13.640 1917.670 13.700 ;
      LAYER met2 ;
        RECT 1890.530 14.010 1890.670 15.300 ;
        RECT 1890.530 13.930 1890.900 14.010 ;
        RECT 1890.530 13.870 1890.960 13.930 ;
        RECT 1890.700 13.610 1890.960 13.870 ;
        RECT 1917.380 13.610 1917.640 13.930 ;
        RECT 1917.440 7.890 1917.580 13.610 ;
        RECT 1917.440 7.750 1918.040 7.890 ;
        RECT 1917.900 2.400 1918.040 7.750 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.090 14.125 1907.230 15.300 ;
        RECT 1907.020 13.755 1907.300 14.125 ;
        RECT 1935.770 13.755 1936.050 14.125 ;
        RECT 1935.840 2.400 1935.980 13.755 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
      LAYER met3 ;
        RECT 1919.430 14.470 1935.370 14.770 ;
        RECT 1906.995 14.090 1907.325 14.105 ;
        RECT 1919.430 14.090 1919.730 14.470 ;
        RECT 1906.995 13.790 1919.730 14.090 ;
        RECT 1935.070 14.090 1935.370 14.470 ;
        RECT 1935.745 14.090 1936.075 14.105 ;
        RECT 1935.070 13.790 1936.075 14.090 ;
        RECT 1906.995 13.775 1907.325 13.790 ;
        RECT 1935.745 13.775 1936.075 13.790 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.650 14.520 1923.790 15.300 ;
        RECT 1923.650 14.380 1924.940 14.520 ;
        RECT 1924.800 14.125 1924.940 14.380 ;
        RECT 1924.730 13.755 1925.010 14.125 ;
        RECT 1952.790 13.330 1953.070 13.445 ;
        RECT 1952.790 13.190 1953.460 13.330 ;
        RECT 1952.790 13.075 1953.070 13.190 ;
        RECT 1953.320 2.400 1953.460 13.190 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER met3 ;
        RECT 1924.705 14.090 1925.035 14.105 ;
        RECT 1924.705 13.790 1934.450 14.090 ;
        RECT 1924.705 13.775 1925.035 13.790 ;
        RECT 1934.150 13.410 1934.450 13.790 ;
        RECT 1952.765 13.410 1953.095 13.425 ;
        RECT 1934.150 13.110 1953.095 13.410 ;
        RECT 1952.765 13.095 1953.095 13.110 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1966.110 14.520 1966.430 14.580 ;
        RECT 1970.250 14.520 1970.570 14.580 ;
        RECT 1966.110 14.380 1970.570 14.520 ;
        RECT 1966.110 14.320 1966.430 14.380 ;
        RECT 1970.250 14.320 1970.570 14.380 ;
      LAYER met2 ;
        RECT 1940.210 14.125 1940.350 15.300 ;
        RECT 1966.140 14.290 1966.400 14.610 ;
        RECT 1970.280 14.520 1970.540 14.610 ;
        RECT 1970.280 14.380 1971.400 14.520 ;
        RECT 1970.280 14.290 1970.540 14.380 ;
        RECT 1966.200 14.125 1966.340 14.290 ;
        RECT 1940.140 13.755 1940.420 14.125 ;
        RECT 1966.130 13.755 1966.410 14.125 ;
        RECT 1971.260 2.400 1971.400 14.380 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
      LAYER met3 ;
        RECT 1940.115 14.090 1940.445 14.105 ;
        RECT 1966.105 14.090 1966.435 14.105 ;
        RECT 1940.115 13.790 1966.435 14.090 ;
        RECT 1940.115 13.775 1940.445 13.790 ;
        RECT 1966.105 13.775 1966.435 13.790 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.770 14.805 1956.910 15.300 ;
        RECT 1956.700 14.435 1956.980 14.805 ;
        RECT 1987.750 13.330 1988.030 13.445 ;
        RECT 1987.750 13.190 1988.880 13.330 ;
        RECT 1987.750 13.075 1988.030 13.190 ;
        RECT 1988.740 2.400 1988.880 13.190 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
      LAYER met3 ;
        RECT 1987.470 16.810 1987.850 16.820 ;
        RECT 1960.830 16.510 1987.850 16.810 ;
        RECT 1956.675 14.770 1957.005 14.785 ;
        RECT 1960.830 14.770 1961.130 16.510 ;
        RECT 1987.470 16.500 1987.850 16.510 ;
        RECT 1956.675 14.470 1961.130 14.770 ;
        RECT 1956.675 14.455 1957.005 14.470 ;
        RECT 1987.725 13.420 1988.055 13.425 ;
        RECT 1987.470 13.410 1988.055 13.420 ;
        RECT 1987.470 13.110 1988.280 13.410 ;
        RECT 1987.470 13.100 1988.055 13.110 ;
        RECT 1987.725 13.095 1988.055 13.100 ;
      LAYER met4 ;
        RECT 1987.495 16.495 1987.825 16.825 ;
        RECT 1987.510 13.425 1987.810 16.495 ;
        RECT 1987.495 13.095 1987.825 13.425 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1973.240 14.520 1973.560 14.580 ;
        RECT 2004.290 14.520 2004.610 14.580 ;
        RECT 1973.240 14.380 2004.610 14.520 ;
        RECT 1973.240 14.320 1973.560 14.380 ;
        RECT 2004.290 14.320 2004.610 14.380 ;
      LAYER met2 ;
        RECT 1973.330 14.610 1973.470 15.300 ;
        RECT 1973.270 14.290 1973.530 14.610 ;
        RECT 2004.320 14.520 2004.580 14.610 ;
        RECT 2004.320 14.380 2005.900 14.520 ;
        RECT 2004.320 14.290 2004.580 14.380 ;
        RECT 2005.760 7.890 2005.900 14.380 ;
        RECT 2005.760 7.750 2006.820 7.890 ;
        RECT 2006.680 2.400 2006.820 7.750 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.890 14.010 1990.030 15.300 ;
        RECT 1989.890 13.870 1990.260 14.010 ;
        RECT 1990.120 6.645 1990.260 13.870 ;
        RECT 1990.050 6.275 1990.330 6.645 ;
        RECT 2024.090 6.275 2024.370 6.645 ;
        RECT 2024.160 2.400 2024.300 6.275 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
      LAYER met3 ;
        RECT 1990.025 6.610 1990.355 6.625 ;
        RECT 2024.065 6.610 2024.395 6.625 ;
        RECT 1990.025 6.310 2024.395 6.610 ;
        RECT 1990.025 6.295 1990.355 6.310 ;
        RECT 2024.065 6.295 2024.395 6.310 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.450 14.010 2006.590 15.300 ;
        RECT 2006.450 13.870 2006.820 14.010 ;
        RECT 2006.680 10.045 2006.820 13.870 ;
        RECT 2006.610 9.675 2006.890 10.045 ;
        RECT 2042.030 9.675 2042.310 10.045 ;
        RECT 2042.100 2.400 2042.240 9.675 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
      LAYER met3 ;
        RECT 2006.585 10.010 2006.915 10.025 ;
        RECT 2042.005 10.010 2042.335 10.025 ;
        RECT 2006.585 9.710 2042.335 10.010 ;
        RECT 2006.585 9.695 2006.915 9.710 ;
        RECT 2042.005 9.695 2042.335 9.710 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.050 14.180 765.370 14.240 ;
        RECT 814.040 14.180 814.360 14.240 ;
        RECT 765.050 14.040 814.360 14.180 ;
        RECT 765.050 13.980 765.370 14.040 ;
        RECT 814.040 13.980 814.360 14.040 ;
      LAYER met2 ;
        RECT 814.130 14.270 814.270 15.300 ;
        RECT 765.080 13.950 765.340 14.270 ;
        RECT 814.070 13.950 814.330 14.270 ;
        RECT 765.140 2.400 765.280 13.950 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2022.920 14.180 2023.240 14.240 ;
        RECT 2058.570 14.180 2058.890 14.240 ;
        RECT 2022.920 14.040 2058.890 14.180 ;
        RECT 2022.920 13.980 2023.240 14.040 ;
        RECT 2058.570 13.980 2058.890 14.040 ;
      LAYER met2 ;
        RECT 2023.010 14.270 2023.150 15.300 ;
        RECT 2022.950 13.950 2023.210 14.270 ;
        RECT 2058.600 13.950 2058.860 14.270 ;
        RECT 2058.660 7.890 2058.800 13.950 ;
        RECT 2058.660 7.750 2059.720 7.890 ;
        RECT 2059.580 2.400 2059.720 7.750 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.570 14.010 2039.710 15.300 ;
        RECT 2039.570 13.870 2039.940 14.010 ;
        RECT 2039.800 0.525 2039.940 13.870 ;
        RECT 2039.730 0.155 2040.010 0.525 ;
        RECT 2076.530 0.410 2076.810 0.525 ;
        RECT 2077.310 0.410 2077.870 2.400 ;
        RECT 2076.530 0.270 2077.870 0.410 ;
        RECT 2076.530 0.155 2076.810 0.270 ;
        RECT 2077.310 -4.800 2077.870 0.270 ;
      LAYER met3 ;
        RECT 2039.705 0.490 2040.035 0.505 ;
        RECT 2076.505 0.490 2076.835 0.505 ;
        RECT 2039.705 0.190 2076.835 0.490 ;
        RECT 2039.705 0.175 2040.035 0.190 ;
        RECT 2076.505 0.175 2076.835 0.190 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2056.130 14.010 2056.270 15.300 ;
        RECT 2055.900 13.870 2056.270 14.010 ;
        RECT 2055.900 3.245 2056.040 13.870 ;
        RECT 2055.830 2.875 2056.110 3.245 ;
        RECT 2094.930 2.875 2095.210 3.245 ;
        RECT 2095.000 2.400 2095.140 2.875 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
      LAYER met3 ;
        RECT 2055.805 3.210 2056.135 3.225 ;
        RECT 2094.905 3.210 2095.235 3.225 ;
        RECT 2055.805 2.910 2095.235 3.210 ;
        RECT 2055.805 2.895 2056.135 2.910 ;
        RECT 2094.905 2.895 2095.235 2.910 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.690 14.010 2072.830 15.300 ;
        RECT 2072.690 13.870 2073.060 14.010 ;
        RECT 2072.920 2.565 2073.060 13.870 ;
        RECT 2072.850 2.195 2073.130 2.565 ;
        RECT 2112.730 1.770 2113.290 2.400 ;
        RECT 2113.790 1.770 2114.070 1.885 ;
        RECT 2112.730 1.630 2114.070 1.770 ;
        RECT 2112.730 -4.800 2113.290 1.630 ;
        RECT 2113.790 1.515 2114.070 1.630 ;
      LAYER met3 ;
        RECT 2072.825 2.530 2073.155 2.545 ;
        RECT 2072.825 2.230 2111.550 2.530 ;
        RECT 2072.825 2.215 2073.155 2.230 ;
        RECT 2111.250 1.850 2111.550 2.230 ;
        RECT 2113.765 1.850 2114.095 1.865 ;
        RECT 2111.250 1.550 2114.095 1.850 ;
        RECT 2113.765 1.535 2114.095 1.550 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.250 14.010 2089.390 15.300 ;
        RECT 2089.250 13.870 2089.620 14.010 ;
        RECT 2089.480 3.925 2089.620 13.870 ;
        RECT 2089.410 3.555 2089.690 3.925 ;
        RECT 2130.810 3.555 2131.090 3.925 ;
        RECT 2130.880 2.400 2131.020 3.555 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
      LAYER met3 ;
        RECT 2089.385 3.890 2089.715 3.905 ;
        RECT 2130.785 3.890 2131.115 3.905 ;
        RECT 2089.385 3.590 2131.115 3.890 ;
        RECT 2089.385 3.575 2089.715 3.590 ;
        RECT 2130.785 3.575 2131.115 3.590 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.810 14.805 2105.950 15.300 ;
        RECT 2105.740 14.435 2106.020 14.805 ;
        RECT 2145.990 13.075 2146.270 13.445 ;
        RECT 2146.060 1.770 2146.200 13.075 ;
        RECT 2148.150 1.770 2148.710 2.400 ;
        RECT 2146.060 1.630 2148.710 1.770 ;
        RECT 2148.150 -4.800 2148.710 1.630 ;
      LAYER met3 ;
        RECT 2105.715 14.770 2106.045 14.785 ;
        RECT 2105.715 14.470 2146.050 14.770 ;
        RECT 2105.715 14.455 2106.045 14.470 ;
        RECT 2145.750 13.425 2146.050 14.470 ;
        RECT 2145.750 13.110 2146.295 13.425 ;
        RECT 2145.965 13.095 2146.295 13.110 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.370 14.010 2122.510 15.300 ;
        RECT 2122.370 13.870 2122.740 14.010 ;
        RECT 2122.600 10.725 2122.740 13.870 ;
        RECT 2122.530 10.355 2122.810 10.725 ;
        RECT 2166.230 10.355 2166.510 10.725 ;
        RECT 2166.300 2.400 2166.440 10.355 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
      LAYER met3 ;
        RECT 2122.505 10.690 2122.835 10.705 ;
        RECT 2166.205 10.690 2166.535 10.705 ;
        RECT 2122.505 10.390 2166.535 10.690 ;
        RECT 2122.505 10.375 2122.835 10.390 ;
        RECT 2166.205 10.375 2166.535 10.390 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.930 14.010 2139.070 15.300 ;
        RECT 2138.700 13.870 2139.070 14.010 ;
        RECT 2138.700 10.045 2138.840 13.870 ;
        RECT 2138.630 9.675 2138.910 10.045 ;
        RECT 2183.710 9.675 2183.990 10.045 ;
        RECT 2183.780 2.400 2183.920 9.675 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
      LAYER met3 ;
        RECT 2138.605 10.010 2138.935 10.025 ;
        RECT 2183.685 10.010 2184.015 10.025 ;
        RECT 2138.605 9.710 2184.015 10.010 ;
        RECT 2138.605 9.695 2138.935 9.710 ;
        RECT 2183.685 9.695 2184.015 9.710 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2155.630 6.700 2155.950 6.760 ;
        RECT 2199.790 6.700 2200.110 6.760 ;
        RECT 2155.630 6.560 2200.110 6.700 ;
        RECT 2155.630 6.500 2155.950 6.560 ;
        RECT 2199.790 6.500 2200.110 6.560 ;
      LAYER met2 ;
        RECT 2155.490 14.010 2155.630 15.300 ;
        RECT 2155.490 13.870 2155.860 14.010 ;
        RECT 2155.720 6.790 2155.860 13.870 ;
        RECT 2155.660 6.470 2155.920 6.790 ;
        RECT 2199.820 6.470 2200.080 6.790 ;
        RECT 2199.880 1.090 2200.020 6.470 ;
        RECT 2201.510 1.090 2202.070 2.400 ;
        RECT 2199.880 0.950 2202.070 1.090 ;
        RECT 2201.510 -4.800 2202.070 0.950 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.050 14.010 2172.190 15.300 ;
        RECT 2172.050 13.870 2172.420 14.010 ;
        RECT 2172.280 8.685 2172.420 13.870 ;
        RECT 2172.210 8.315 2172.490 8.685 ;
        RECT 2219.130 8.315 2219.410 8.685 ;
        RECT 2219.200 2.400 2219.340 8.315 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
      LAYER met3 ;
        RECT 2172.185 8.650 2172.515 8.665 ;
        RECT 2219.105 8.650 2219.435 8.665 ;
        RECT 2172.185 8.350 2219.435 8.650 ;
        RECT 2172.185 8.335 2172.515 8.350 ;
        RECT 2219.105 8.335 2219.435 8.350 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.690 14.010 830.830 15.300 ;
        RECT 830.460 13.870 830.830 14.010 ;
        RECT 830.460 12.085 830.600 13.870 ;
        RECT 783.010 11.715 783.290 12.085 ;
        RECT 830.390 11.715 830.670 12.085 ;
        RECT 783.080 2.400 783.220 11.715 ;
        RECT 782.870 -4.800 783.430 2.400 ;
      LAYER met3 ;
        RECT 782.985 12.050 783.315 12.065 ;
        RECT 830.365 12.050 830.695 12.065 ;
        RECT 782.985 11.750 830.695 12.050 ;
        RECT 782.985 11.735 783.315 11.750 ;
        RECT 830.365 11.735 830.695 11.750 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.610 14.010 2188.750 15.300 ;
        RECT 2188.610 13.870 2188.980 14.010 ;
        RECT 2188.840 10.045 2188.980 13.870 ;
        RECT 2188.770 9.675 2189.050 10.045 ;
        RECT 2237.070 9.675 2237.350 10.045 ;
        RECT 2237.140 2.400 2237.280 9.675 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
      LAYER met3 ;
        RECT 2188.745 10.010 2189.075 10.025 ;
        RECT 2237.045 10.010 2237.375 10.025 ;
        RECT 2188.745 9.710 2237.375 10.010 ;
        RECT 2188.745 9.695 2189.075 9.710 ;
        RECT 2237.045 9.695 2237.375 9.710 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.170 14.010 2205.310 15.300 ;
        RECT 2205.170 13.870 2205.540 14.010 ;
        RECT 2205.400 13.445 2205.540 13.870 ;
        RECT 2205.330 13.075 2205.610 13.445 ;
        RECT 2254.550 13.075 2254.830 13.445 ;
        RECT 2254.620 2.400 2254.760 13.075 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
      LAYER met3 ;
        RECT 2205.305 13.410 2205.635 13.425 ;
        RECT 2254.525 13.410 2254.855 13.425 ;
        RECT 2205.305 13.110 2254.855 13.410 ;
        RECT 2205.305 13.095 2205.635 13.110 ;
        RECT 2254.525 13.095 2254.855 13.110 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2221.410 0.580 2221.730 0.640 ;
        RECT 2270.630 0.580 2270.950 0.640 ;
        RECT 2221.410 0.440 2270.950 0.580 ;
        RECT 2221.410 0.380 2221.730 0.440 ;
        RECT 2270.630 0.380 2270.950 0.440 ;
      LAYER met2 ;
        RECT 2221.730 14.010 2221.870 15.300 ;
        RECT 2221.500 13.870 2221.870 14.010 ;
        RECT 2221.500 0.670 2221.640 13.870 ;
        RECT 2221.440 0.350 2221.700 0.670 ;
        RECT 2270.660 0.410 2270.920 0.670 ;
        RECT 2272.350 0.410 2272.910 2.400 ;
        RECT 2270.660 0.350 2272.910 0.410 ;
        RECT 2270.720 0.270 2272.910 0.350 ;
        RECT 2272.350 -4.800 2272.910 0.270 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.290 14.010 2238.430 15.300 ;
        RECT 2238.290 13.870 2238.660 14.010 ;
        RECT 2238.520 2.565 2238.660 13.870 ;
        RECT 2289.580 2.990 2290.640 3.130 ;
        RECT 2238.450 2.195 2238.730 2.565 ;
        RECT 2288.590 2.450 2288.870 2.565 ;
        RECT 2289.580 2.450 2289.720 2.990 ;
        RECT 2288.590 2.310 2289.720 2.450 ;
        RECT 2290.500 2.400 2290.640 2.990 ;
        RECT 2288.590 2.195 2288.870 2.310 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
      LAYER met3 ;
        RECT 2238.425 2.530 2238.755 2.545 ;
        RECT 2288.565 2.530 2288.895 2.545 ;
        RECT 2238.425 2.230 2288.895 2.530 ;
        RECT 2238.425 2.215 2238.755 2.230 ;
        RECT 2288.565 2.215 2288.895 2.230 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2254.990 6.700 2255.310 6.760 ;
        RECT 2306.510 6.700 2306.830 6.760 ;
        RECT 2254.990 6.560 2306.830 6.700 ;
        RECT 2254.990 6.500 2255.310 6.560 ;
        RECT 2306.510 6.500 2306.830 6.560 ;
      LAYER met2 ;
        RECT 2254.850 14.010 2254.990 15.300 ;
        RECT 2254.850 13.870 2255.220 14.010 ;
        RECT 2255.080 6.790 2255.220 13.870 ;
        RECT 2255.020 6.470 2255.280 6.790 ;
        RECT 2306.540 6.470 2306.800 6.790 ;
        RECT 2306.600 3.810 2306.740 6.470 ;
        RECT 2306.600 3.670 2308.120 3.810 ;
        RECT 2307.980 2.400 2308.120 3.670 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2271.550 6.360 2271.870 6.420 ;
        RECT 2325.370 6.360 2325.690 6.420 ;
        RECT 2271.550 6.220 2325.690 6.360 ;
        RECT 2271.550 6.160 2271.870 6.220 ;
        RECT 2325.370 6.160 2325.690 6.220 ;
      LAYER met2 ;
        RECT 2271.410 14.010 2271.550 15.300 ;
        RECT 2271.410 13.870 2271.780 14.010 ;
        RECT 2271.640 6.450 2271.780 13.870 ;
        RECT 2271.580 6.130 2271.840 6.450 ;
        RECT 2325.400 6.360 2325.660 6.450 ;
        RECT 2325.400 6.220 2326.060 6.360 ;
        RECT 2325.400 6.130 2325.660 6.220 ;
        RECT 2325.920 2.400 2326.060 6.220 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.970 13.870 2288.110 15.300 ;
        RECT 2287.970 13.730 2288.340 13.870 ;
        RECT 2288.200 0.525 2288.340 13.730 ;
        RECT 2342.480 2.990 2343.540 3.130 ;
        RECT 2342.480 0.525 2342.620 2.990 ;
        RECT 2343.400 2.400 2343.540 2.990 ;
        RECT 2288.130 0.155 2288.410 0.525 ;
        RECT 2342.410 0.155 2342.690 0.525 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
      LAYER met3 ;
        RECT 2288.105 0.490 2288.435 0.505 ;
        RECT 2342.385 0.490 2342.715 0.505 ;
        RECT 2288.105 0.190 2342.715 0.490 ;
        RECT 2288.105 0.175 2288.435 0.190 ;
        RECT 2342.385 0.175 2342.715 0.190 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2304.210 0.580 2304.530 0.640 ;
        RECT 2362.170 0.580 2362.490 0.640 ;
        RECT 2304.210 0.440 2362.490 0.580 ;
        RECT 2304.210 0.380 2304.530 0.440 ;
        RECT 2362.170 0.380 2362.490 0.440 ;
      LAYER met2 ;
        RECT 2304.530 13.870 2304.670 15.300 ;
        RECT 2304.300 13.730 2304.670 13.870 ;
        RECT 2304.300 0.670 2304.440 13.730 ;
        RECT 2304.240 0.350 2304.500 0.670 ;
        RECT 2361.130 0.410 2361.690 2.400 ;
        RECT 2362.200 0.410 2362.460 0.670 ;
        RECT 2361.130 0.350 2362.460 0.410 ;
        RECT 2361.130 0.270 2362.400 0.350 ;
        RECT 2361.130 -4.800 2361.690 0.270 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.090 14.805 2321.230 15.300 ;
        RECT 2321.020 14.435 2321.300 14.805 ;
        RECT 2376.910 13.330 2377.190 13.445 ;
        RECT 2376.910 13.190 2378.960 13.330 ;
        RECT 2376.910 13.075 2377.190 13.190 ;
        RECT 2378.820 2.400 2378.960 13.190 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
      LAYER met3 ;
        RECT 2335.270 15.150 2353.050 15.450 ;
        RECT 2320.995 14.770 2321.325 14.785 ;
        RECT 2335.270 14.770 2335.570 15.150 ;
        RECT 2320.995 14.470 2335.570 14.770 ;
        RECT 2320.995 14.455 2321.325 14.470 ;
        RECT 2352.750 14.090 2353.050 15.150 ;
        RECT 2352.750 13.790 2354.890 14.090 ;
        RECT 2354.590 13.410 2354.890 13.790 ;
        RECT 2376.885 13.410 2377.215 13.425 ;
        RECT 2354.590 13.110 2377.215 13.410 ;
        RECT 2376.885 13.095 2377.215 13.110 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2337.790 6.700 2338.110 6.760 ;
        RECT 2364.930 6.700 2365.250 6.760 ;
        RECT 2337.790 6.560 2365.250 6.700 ;
        RECT 2337.790 6.500 2338.110 6.560 ;
        RECT 2364.930 6.500 2365.250 6.560 ;
        RECT 2364.930 5.680 2365.250 5.740 ;
        RECT 2394.370 5.680 2394.690 5.740 ;
        RECT 2364.930 5.540 2394.690 5.680 ;
        RECT 2364.930 5.480 2365.250 5.540 ;
        RECT 2394.370 5.480 2394.690 5.540 ;
      LAYER met2 ;
        RECT 2337.650 14.010 2337.790 15.300 ;
        RECT 2337.650 13.870 2338.020 14.010 ;
        RECT 2337.880 6.790 2338.020 13.870 ;
        RECT 2337.820 6.470 2338.080 6.790 ;
        RECT 2364.960 6.470 2365.220 6.790 ;
        RECT 2365.020 5.770 2365.160 6.470 ;
        RECT 2394.460 5.770 2395.060 5.850 ;
        RECT 2364.960 5.450 2365.220 5.770 ;
        RECT 2394.400 5.710 2395.060 5.770 ;
        RECT 2394.400 5.450 2394.660 5.710 ;
        RECT 2394.920 1.770 2395.060 5.710 ;
        RECT 2396.550 1.770 2397.110 2.400 ;
        RECT 2394.920 1.630 2397.110 1.770 ;
        RECT 2396.550 -4.800 2397.110 1.630 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.250 14.010 847.390 15.300 ;
        RECT 847.020 13.870 847.390 14.010 ;
        RECT 800.560 2.990 801.620 3.130 ;
        RECT 800.560 2.400 800.700 2.990 ;
        RECT 801.480 2.565 801.620 2.990 ;
        RECT 847.020 2.565 847.160 13.870 ;
        RECT 800.350 -4.800 800.910 2.400 ;
        RECT 801.410 2.195 801.690 2.565 ;
        RECT 846.950 2.195 847.230 2.565 ;
      LAYER met3 ;
        RECT 801.385 2.530 801.715 2.545 ;
        RECT 846.925 2.530 847.255 2.545 ;
        RECT 801.385 2.230 847.255 2.530 ;
        RECT 801.385 2.215 801.715 2.230 ;
        RECT 846.925 2.215 847.255 2.230 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2806.990 0.580 2807.310 0.640 ;
        RECT 2905.890 0.580 2906.210 0.640 ;
        RECT 2806.990 0.440 2906.210 0.580 ;
        RECT 2806.990 0.380 2807.310 0.440 ;
        RECT 2905.890 0.380 2906.210 0.440 ;
      LAYER met2 ;
        RECT 2806.850 14.010 2806.990 15.300 ;
        RECT 2806.850 13.870 2807.220 14.010 ;
        RECT 2807.080 0.670 2807.220 13.870 ;
        RECT 2807.020 0.350 2807.280 0.670 ;
        RECT 2904.850 0.410 2905.410 2.400 ;
        RECT 2905.920 0.410 2906.180 0.670 ;
        RECT 2904.850 0.350 2906.180 0.410 ;
        RECT 2904.850 0.270 2906.120 0.350 ;
        RECT 2904.850 -4.800 2905.410 0.270 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2812.370 14.010 2812.510 15.300 ;
        RECT 2812.370 13.870 2812.740 14.010 ;
        RECT 2812.600 1.205 2812.740 13.870 ;
        RECT 2812.530 0.835 2812.810 1.205 ;
        RECT 2909.130 1.090 2909.410 1.205 ;
        RECT 2910.830 1.090 2911.390 2.400 ;
        RECT 2909.130 0.950 2911.390 1.090 ;
        RECT 2909.130 0.835 2909.410 0.950 ;
        RECT 2910.830 -4.800 2911.390 0.950 ;
      LAYER met3 ;
        RECT 2812.505 1.170 2812.835 1.185 ;
        RECT 2909.105 1.170 2909.435 1.185 ;
        RECT 2812.505 0.870 2909.435 1.170 ;
        RECT 2812.505 0.855 2812.835 0.870 ;
        RECT 2909.105 0.855 2909.435 0.870 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2817.890 14.010 2818.030 15.300 ;
        RECT 2817.890 13.870 2818.260 14.010 ;
        RECT 2818.120 0.525 2818.260 13.870 ;
        RECT 2818.050 0.155 2818.330 0.525 ;
        RECT 2916.810 0.410 2917.370 2.400 ;
        RECT 2917.870 0.410 2918.150 0.525 ;
        RECT 2916.810 0.270 2918.150 0.410 ;
        RECT 2916.810 -4.800 2917.370 0.270 ;
        RECT 2917.870 0.155 2918.150 0.270 ;
      LAYER met3 ;
        RECT 2818.025 0.490 2818.355 0.505 ;
        RECT 2917.845 0.490 2918.175 0.505 ;
        RECT 2818.025 0.190 2918.175 0.490 ;
        RECT 2818.025 0.175 2818.355 0.190 ;
        RECT 2917.845 0.175 2918.175 0.190 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
        RECT 81.040 1634.330 82.640 1637.430 ;
        RECT 81.040 1454.330 82.640 1457.430 ;
        RECT 81.040 1274.330 82.640 1277.430 ;
        RECT 81.040 1094.330 82.640 1097.430 ;
        RECT 81.040 914.330 82.640 917.430 ;
        RECT 81.040 734.330 82.640 737.430 ;
        RECT 81.040 554.330 82.640 557.430 ;
        RECT 81.040 374.330 82.640 377.430 ;
        RECT 81.040 194.330 82.640 197.430 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
        RECT 234.640 1634.330 236.240 1637.430 ;
        RECT 234.640 1454.330 236.240 1457.430 ;
        RECT 234.640 1274.330 236.240 1277.430 ;
        RECT 234.640 1094.330 236.240 1097.430 ;
        RECT 234.640 914.330 236.240 917.430 ;
        RECT 234.640 734.330 236.240 737.430 ;
        RECT 234.640 554.330 236.240 557.430 ;
        RECT 234.640 374.330 236.240 377.430 ;
        RECT 234.640 194.330 236.240 197.430 ;
        RECT 368.970 -38.270 372.070 3557.950 ;
        RECT 388.240 1634.330 389.840 1637.430 ;
        RECT 541.840 1634.330 543.440 1637.430 ;
        RECT 388.240 1454.330 389.840 1457.430 ;
        RECT 541.840 1454.330 543.440 1457.430 ;
        RECT 388.240 1274.330 389.840 1277.430 ;
        RECT 541.840 1274.330 543.440 1277.430 ;
        RECT 388.240 1094.330 389.840 1097.430 ;
        RECT 541.840 1094.330 543.440 1097.430 ;
        RECT 388.240 914.330 389.840 917.430 ;
        RECT 541.840 914.330 543.440 917.430 ;
        RECT 388.240 734.330 389.840 737.430 ;
        RECT 541.840 734.330 543.440 737.430 ;
        RECT 388.240 554.330 389.840 557.430 ;
        RECT 541.840 554.330 543.440 557.430 ;
        RECT 388.240 374.330 389.840 377.430 ;
        RECT 541.840 374.330 543.440 377.430 ;
        RECT 388.240 194.330 389.840 197.430 ;
        RECT 541.840 194.330 543.440 197.430 ;
        RECT 548.970 -38.270 552.070 3557.950 ;
        RECT 695.440 1634.330 697.040 1637.430 ;
        RECT 695.440 1454.330 697.040 1457.430 ;
        RECT 695.440 1274.330 697.040 1277.430 ;
        RECT 695.440 1094.330 697.040 1097.430 ;
        RECT 695.440 914.330 697.040 917.430 ;
        RECT 695.440 734.330 697.040 737.430 ;
        RECT 695.440 554.330 697.040 557.430 ;
        RECT 695.440 374.330 697.040 377.430 ;
        RECT 695.440 194.330 697.040 197.430 ;
        RECT 728.970 -38.270 732.070 3557.950 ;
        RECT 849.040 1634.330 850.640 1637.430 ;
        RECT 849.040 1454.330 850.640 1457.430 ;
        RECT 849.040 1274.330 850.640 1277.430 ;
        RECT 849.040 1094.330 850.640 1097.430 ;
        RECT 849.040 914.330 850.640 917.430 ;
        RECT 849.040 734.330 850.640 737.430 ;
        RECT 849.040 554.330 850.640 557.430 ;
        RECT 849.040 374.330 850.640 377.430 ;
        RECT 849.040 194.330 850.640 197.430 ;
        RECT 908.970 -38.270 912.070 3557.950 ;
        RECT 1002.640 1634.330 1004.240 1637.430 ;
        RECT 1002.640 1454.330 1004.240 1457.430 ;
        RECT 1002.640 1274.330 1004.240 1277.430 ;
        RECT 1002.640 1094.330 1004.240 1097.430 ;
        RECT 1002.640 914.330 1004.240 917.430 ;
        RECT 1002.640 734.330 1004.240 737.430 ;
        RECT 1002.640 554.330 1004.240 557.430 ;
        RECT 1002.640 374.330 1004.240 377.430 ;
        RECT 1002.640 194.330 1004.240 197.430 ;
        RECT 1088.970 -38.270 1092.070 3557.950 ;
        RECT 1156.240 1634.330 1157.840 1637.430 ;
        RECT 1156.240 1454.330 1157.840 1457.430 ;
        RECT 1156.240 1274.330 1157.840 1277.430 ;
        RECT 1156.240 1094.330 1157.840 1097.430 ;
        RECT 1156.240 914.330 1157.840 917.430 ;
        RECT 1156.240 734.330 1157.840 737.430 ;
        RECT 1156.240 554.330 1157.840 557.430 ;
        RECT 1156.240 374.330 1157.840 377.430 ;
        RECT 1156.240 194.330 1157.840 197.430 ;
        RECT 1268.970 -38.270 1272.070 3557.950 ;
        RECT 1309.840 1634.330 1311.440 1637.430 ;
        RECT 1309.840 1454.330 1311.440 1457.430 ;
        RECT 1309.840 1274.330 1311.440 1277.430 ;
        RECT 1309.840 1094.330 1311.440 1097.430 ;
        RECT 1309.840 914.330 1311.440 917.430 ;
        RECT 1309.840 734.330 1311.440 737.430 ;
        RECT 1309.840 554.330 1311.440 557.430 ;
        RECT 1309.840 374.330 1311.440 377.430 ;
        RECT 1309.840 194.330 1311.440 197.430 ;
        RECT 1448.970 -38.270 1452.070 3557.950 ;
        RECT 1463.440 1634.330 1465.040 1637.430 ;
        RECT 1617.040 1634.330 1618.640 1637.430 ;
        RECT 1463.440 1454.330 1465.040 1457.430 ;
        RECT 1617.040 1454.330 1618.640 1457.430 ;
        RECT 1463.440 1274.330 1465.040 1277.430 ;
        RECT 1617.040 1274.330 1618.640 1277.430 ;
        RECT 1463.440 1094.330 1465.040 1097.430 ;
        RECT 1617.040 1094.330 1618.640 1097.430 ;
        RECT 1463.440 914.330 1465.040 917.430 ;
        RECT 1617.040 914.330 1618.640 917.430 ;
        RECT 1463.440 734.330 1465.040 737.430 ;
        RECT 1617.040 734.330 1618.640 737.430 ;
        RECT 1463.440 554.330 1465.040 557.430 ;
        RECT 1617.040 554.330 1618.640 557.430 ;
        RECT 1463.440 374.330 1465.040 377.430 ;
        RECT 1617.040 374.330 1618.640 377.430 ;
        RECT 1463.440 194.330 1465.040 197.430 ;
        RECT 1617.040 194.330 1618.640 197.430 ;
        RECT 1628.970 -38.270 1632.070 3557.950 ;
        RECT 1770.640 1634.330 1772.240 1637.430 ;
        RECT 1770.640 1454.330 1772.240 1457.430 ;
        RECT 1770.640 1274.330 1772.240 1277.430 ;
        RECT 1770.640 1094.330 1772.240 1097.430 ;
        RECT 1770.640 914.330 1772.240 917.430 ;
        RECT 1770.640 734.330 1772.240 737.430 ;
        RECT 1770.640 554.330 1772.240 557.430 ;
        RECT 1770.640 374.330 1772.240 377.430 ;
        RECT 1770.640 194.330 1772.240 197.430 ;
        RECT 1808.970 -38.270 1812.070 3557.950 ;
        RECT 1924.240 1634.330 1925.840 1637.430 ;
        RECT 1924.240 1454.330 1925.840 1457.430 ;
        RECT 1924.240 1274.330 1925.840 1277.430 ;
        RECT 1924.240 1094.330 1925.840 1097.430 ;
        RECT 1924.240 914.330 1925.840 917.430 ;
        RECT 1924.240 734.330 1925.840 737.430 ;
        RECT 1924.240 554.330 1925.840 557.430 ;
        RECT 1924.240 374.330 1925.840 377.430 ;
        RECT 1924.240 194.330 1925.840 197.430 ;
        RECT 1988.970 -38.270 1992.070 3557.950 ;
        RECT 2077.840 1634.330 2079.440 1637.430 ;
        RECT 2077.840 1454.330 2079.440 1457.430 ;
        RECT 2077.840 1274.330 2079.440 1277.430 ;
        RECT 2077.840 1094.330 2079.440 1097.430 ;
        RECT 2077.840 914.330 2079.440 917.430 ;
        RECT 2077.840 734.330 2079.440 737.430 ;
        RECT 2077.840 554.330 2079.440 557.430 ;
        RECT 2077.840 374.330 2079.440 377.430 ;
        RECT 2077.840 194.330 2079.440 197.430 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
        RECT 2231.440 1634.330 2233.040 1637.430 ;
        RECT 2231.440 1454.330 2233.040 1457.430 ;
        RECT 2231.440 1274.330 2233.040 1277.430 ;
        RECT 2231.440 1094.330 2233.040 1097.430 ;
        RECT 2231.440 914.330 2233.040 917.430 ;
        RECT 2231.440 734.330 2233.040 737.430 ;
        RECT 2231.440 554.330 2233.040 557.430 ;
        RECT 2231.440 374.330 2233.040 377.430 ;
        RECT 2231.440 194.330 2233.040 197.430 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
        RECT 2385.040 1634.330 2386.640 1637.430 ;
        RECT 2385.040 1454.330 2386.640 1457.430 ;
        RECT 2385.040 1274.330 2386.640 1277.430 ;
        RECT 2385.040 1094.330 2386.640 1097.430 ;
        RECT 2385.040 914.330 2386.640 917.430 ;
        RECT 2385.040 734.330 2386.640 737.430 ;
        RECT 2385.040 554.330 2386.640 557.430 ;
        RECT 2385.040 374.330 2386.640 377.430 ;
        RECT 2385.040 194.330 2386.640 197.430 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
        RECT 2538.640 1634.330 2540.240 1637.430 ;
        RECT 2692.240 1634.330 2693.840 1637.430 ;
        RECT 2538.640 1454.330 2540.240 1457.430 ;
        RECT 2692.240 1454.330 2693.840 1457.430 ;
        RECT 2538.640 1274.330 2540.240 1277.430 ;
        RECT 2692.240 1274.330 2693.840 1277.430 ;
        RECT 2538.640 1094.330 2540.240 1097.430 ;
        RECT 2692.240 1094.330 2693.840 1097.430 ;
        RECT 2538.640 914.330 2540.240 917.430 ;
        RECT 2692.240 914.330 2693.840 917.430 ;
        RECT 2538.640 734.330 2540.240 737.430 ;
        RECT 2692.240 734.330 2693.840 737.430 ;
        RECT 2538.640 554.330 2540.240 557.430 ;
        RECT 2692.240 554.330 2693.840 557.430 ;
        RECT 2538.640 374.330 2540.240 377.430 ;
        RECT 2692.240 374.330 2693.840 377.430 ;
        RECT 2538.640 194.330 2540.240 197.430 ;
        RECT 2692.240 194.330 2693.840 197.430 ;
        RECT 2708.970 -38.270 2712.070 3557.950 ;
        RECT 2845.840 1634.330 2847.440 1637.430 ;
        RECT 2845.840 1454.330 2847.440 1457.430 ;
        RECT 2845.840 1274.330 2847.440 1277.430 ;
        RECT 2845.840 1094.330 2847.440 1097.430 ;
        RECT 2845.840 914.330 2847.440 917.430 ;
        RECT 2845.840 734.330 2847.440 737.430 ;
        RECT 2845.840 554.330 2847.440 557.430 ;
        RECT 2845.840 374.330 2847.440 377.430 ;
        RECT 2845.840 194.330 2847.440 197.430 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
        RECT -43.630 914.330 2963.250 917.430 ;
        RECT -43.630 734.330 2963.250 737.430 ;
        RECT -43.630 554.330 2963.250 557.430 ;
        RECT -43.630 374.330 2963.250 377.430 ;
        RECT -43.630 194.330 2963.250 197.430 ;
        RECT -43.630 14.330 2963.250 17.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 46.170 -38.270 49.270 3557.950 ;
        RECT 226.170 -38.270 229.270 3557.950 ;
        RECT 406.170 -38.270 409.270 3557.950 ;
        RECT 586.170 -38.270 589.270 3557.950 ;
        RECT 766.170 -38.270 769.270 3557.950 ;
        RECT 946.170 -38.270 949.270 3557.950 ;
        RECT 1126.170 -38.270 1129.270 3557.950 ;
        RECT 1306.170 1774.900 1309.270 3557.950 ;
        RECT 1486.170 -38.270 1489.270 3557.950 ;
        RECT 1666.170 -38.270 1669.270 3557.950 ;
        RECT 1846.170 1774.900 1849.270 3557.950 ;
        RECT 2026.170 -38.270 2029.270 3557.950 ;
        RECT 2206.170 -38.270 2209.270 3557.950 ;
        RECT 2386.170 1774.900 2389.270 3557.950 ;
        RECT 2566.170 -38.270 2569.270 3557.950 ;
        RECT 2746.170 -38.270 2749.270 3557.950 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -43.630 3471.530 2963.250 3474.630 ;
        RECT -43.630 3291.530 2963.250 3294.630 ;
        RECT -43.630 3111.530 2963.250 3114.630 ;
        RECT -43.630 2931.530 2963.250 2934.630 ;
        RECT -43.630 2751.530 2963.250 2754.630 ;
        RECT -43.630 2571.530 2963.250 2574.630 ;
        RECT -43.630 2391.530 2963.250 2394.630 ;
        RECT -43.630 2211.530 2963.250 2214.630 ;
        RECT -43.630 2031.530 2963.250 2034.630 ;
        RECT -43.630 1851.530 2963.250 1854.630 ;
        RECT -43.630 1671.530 2963.250 1674.630 ;
        RECT -43.630 1491.530 2963.250 1494.630 ;
        RECT -43.630 1311.530 2963.250 1314.630 ;
        RECT -43.630 1131.530 2963.250 1134.630 ;
        RECT -43.630 951.530 2963.250 954.630 ;
        RECT -43.630 771.530 2963.250 774.630 ;
        RECT -43.630 591.530 2963.250 594.630 ;
        RECT -43.630 411.530 2963.250 414.630 ;
        RECT -43.630 231.530 2963.250 234.630 ;
        RECT -43.630 51.530 2963.250 54.630 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 83.370 -38.270 86.470 3557.950 ;
        RECT 263.370 -38.270 266.470 3557.950 ;
        RECT 443.370 -38.270 446.470 3557.950 ;
        RECT 623.370 -38.270 626.470 3557.950 ;
        RECT 803.370 -38.270 806.470 3557.950 ;
        RECT 983.370 -38.270 986.470 3557.950 ;
        RECT 1163.370 -38.270 1166.470 3557.950 ;
        RECT 1343.370 -38.270 1346.470 3557.950 ;
        RECT 1523.370 -38.270 1526.470 3557.950 ;
        RECT 1703.370 -38.270 1706.470 3557.950 ;
        RECT 1883.370 -38.270 1886.470 3557.950 ;
        RECT 2063.370 -38.270 2066.470 3557.950 ;
        RECT 2243.370 -38.270 2246.470 3557.950 ;
        RECT 2423.370 -38.270 2426.470 3557.950 ;
        RECT 2603.370 -38.270 2606.470 3557.950 ;
        RECT 2783.370 -38.270 2786.470 3557.950 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -43.630 3328.730 2963.250 3331.830 ;
        RECT -43.630 3148.730 2963.250 3151.830 ;
        RECT -43.630 2968.730 2963.250 2971.830 ;
        RECT -43.630 2788.730 2963.250 2791.830 ;
        RECT -43.630 2608.730 2963.250 2611.830 ;
        RECT -43.630 2428.730 2963.250 2431.830 ;
        RECT -43.630 2248.730 2963.250 2251.830 ;
        RECT -43.630 2068.730 2963.250 2071.830 ;
        RECT -43.630 1888.730 2963.250 1891.830 ;
        RECT -43.630 1708.730 2963.250 1711.830 ;
        RECT -43.630 1528.730 2963.250 1531.830 ;
        RECT -43.630 1348.730 2963.250 1351.830 ;
        RECT -43.630 1168.730 2963.250 1171.830 ;
        RECT -43.630 988.730 2963.250 991.830 ;
        RECT -43.630 808.730 2963.250 811.830 ;
        RECT -43.630 628.730 2963.250 631.830 ;
        RECT -43.630 448.730 2963.250 451.830 ;
        RECT -43.630 268.730 2963.250 271.830 ;
        RECT -43.630 88.730 2963.250 91.830 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 120.570 -38.270 123.670 3557.950 ;
        RECT 300.570 -38.270 303.670 3557.950 ;
        RECT 480.570 -38.270 483.670 3557.950 ;
        RECT 660.570 -38.270 663.670 3557.950 ;
        RECT 840.570 -38.270 843.670 3557.950 ;
        RECT 1020.570 -38.270 1023.670 3557.950 ;
        RECT 1200.570 -38.270 1203.670 3557.950 ;
        RECT 1380.570 -38.270 1383.670 3557.950 ;
        RECT 1560.570 -38.270 1563.670 3557.950 ;
        RECT 1740.570 -38.270 1743.670 3557.950 ;
        RECT 1920.570 1774.900 1923.670 3557.950 ;
        RECT 2100.570 -38.270 2103.670 3557.950 ;
        RECT 2280.570 -38.270 2283.670 3557.950 ;
        RECT 2460.570 1774.900 2463.670 3557.950 ;
        RECT 2640.570 -38.270 2643.670 3557.950 ;
        RECT 2820.570 -38.270 2823.670 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3365.930 2963.250 3369.030 ;
        RECT -43.630 3185.930 2963.250 3189.030 ;
        RECT -43.630 3005.930 2963.250 3009.030 ;
        RECT -43.630 2825.930 2963.250 2829.030 ;
        RECT -43.630 2645.930 2963.250 2649.030 ;
        RECT -43.630 2465.930 2963.250 2469.030 ;
        RECT -43.630 2285.930 2963.250 2289.030 ;
        RECT -43.630 2105.930 2963.250 2109.030 ;
        RECT -43.630 1925.930 2963.250 1929.030 ;
        RECT -43.630 1745.930 2963.250 1749.030 ;
        RECT -43.630 1565.930 2963.250 1569.030 ;
        RECT -43.630 1385.930 2963.250 1389.030 ;
        RECT -43.630 1205.930 2963.250 1209.030 ;
        RECT -43.630 1025.930 2963.250 1029.030 ;
        RECT -43.630 845.930 2963.250 849.030 ;
        RECT -43.630 665.930 2963.250 669.030 ;
        RECT -43.630 485.930 2963.250 489.030 ;
        RECT -43.630 305.930 2963.250 309.030 ;
        RECT -43.630 125.930 2963.250 129.030 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 101.970 -38.270 105.070 3557.950 ;
        RECT 281.970 -38.270 285.070 3557.950 ;
        RECT 461.970 1774.900 465.070 3557.950 ;
        RECT 641.970 -38.270 645.070 3557.950 ;
        RECT 821.970 -38.270 825.070 3557.950 ;
        RECT 1001.970 1774.900 1005.070 3557.950 ;
        RECT 1181.970 -38.270 1185.070 3557.950 ;
        RECT 1361.970 -38.270 1365.070 3557.950 ;
        RECT 1541.970 1774.900 1545.070 3557.950 ;
        RECT 1721.970 -38.270 1725.070 3557.950 ;
        RECT 1901.970 -38.270 1905.070 3557.950 ;
        RECT 2081.970 -38.270 2085.070 3557.950 ;
        RECT 2261.970 -38.270 2265.070 3557.950 ;
        RECT 2441.970 -38.270 2445.070 3557.950 ;
        RECT 2621.970 -38.270 2625.070 3557.950 ;
        RECT 2801.970 -38.270 2805.070 3557.950 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -43.630 3347.330 2963.250 3350.430 ;
        RECT -43.630 3167.330 2963.250 3170.430 ;
        RECT -43.630 2987.330 2963.250 2990.430 ;
        RECT -43.630 2807.330 2963.250 2810.430 ;
        RECT -43.630 2627.330 2963.250 2630.430 ;
        RECT -43.630 2447.330 2963.250 2450.430 ;
        RECT -43.630 2267.330 2963.250 2270.430 ;
        RECT -43.630 2087.330 2963.250 2090.430 ;
        RECT -43.630 1907.330 2963.250 1910.430 ;
        RECT -43.630 1727.330 2963.250 1730.430 ;
        RECT -43.630 1547.330 2963.250 1550.430 ;
        RECT -43.630 1367.330 2963.250 1370.430 ;
        RECT -43.630 1187.330 2963.250 1190.430 ;
        RECT -43.630 1007.330 2963.250 1010.430 ;
        RECT -43.630 827.330 2963.250 830.430 ;
        RECT -43.630 647.330 2963.250 650.430 ;
        RECT -43.630 467.330 2963.250 470.430 ;
        RECT -43.630 287.330 2963.250 290.430 ;
        RECT -43.630 107.330 2963.250 110.430 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 139.170 -38.270 142.270 3557.950 ;
        RECT 319.170 -38.270 322.270 3557.950 ;
        RECT 499.170 -38.270 502.270 3557.950 ;
        RECT 679.170 -38.270 682.270 3557.950 ;
        RECT 859.170 -38.270 862.270 3557.950 ;
        RECT 1039.170 -38.270 1042.270 3557.950 ;
        RECT 1219.170 -38.270 1222.270 3557.950 ;
        RECT 1399.170 -38.270 1402.270 3557.950 ;
        RECT 1579.170 -38.270 1582.270 3557.950 ;
        RECT 1759.170 -38.270 1762.270 3557.950 ;
        RECT 1939.170 -38.270 1942.270 3557.950 ;
        RECT 2119.170 -38.270 2122.270 3557.950 ;
        RECT 2299.170 -38.270 2302.270 3557.950 ;
        RECT 2479.170 -38.270 2482.270 3557.950 ;
        RECT 2659.170 -38.270 2662.270 3557.950 ;
        RECT 2839.170 -38.270 2842.270 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3384.530 2963.250 3387.630 ;
        RECT -43.630 3204.530 2963.250 3207.630 ;
        RECT -43.630 3024.530 2963.250 3027.630 ;
        RECT -43.630 2844.530 2963.250 2847.630 ;
        RECT -43.630 2664.530 2963.250 2667.630 ;
        RECT -43.630 2484.530 2963.250 2487.630 ;
        RECT -43.630 2304.530 2963.250 2307.630 ;
        RECT -43.630 2124.530 2963.250 2127.630 ;
        RECT -43.630 1944.530 2963.250 1947.630 ;
        RECT -43.630 1764.530 2963.250 1767.630 ;
        RECT -43.630 1584.530 2963.250 1587.630 ;
        RECT -43.630 1404.530 2963.250 1407.630 ;
        RECT -43.630 1224.530 2963.250 1227.630 ;
        RECT -43.630 1044.530 2963.250 1047.630 ;
        RECT -43.630 864.530 2963.250 867.630 ;
        RECT -43.630 684.530 2963.250 687.630 ;
        RECT -43.630 504.530 2963.250 507.630 ;
        RECT -43.630 324.530 2963.250 327.630 ;
        RECT -43.630 144.530 2963.250 147.630 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 27.570 -38.270 30.670 3557.950 ;
        RECT 157.840 1652.930 159.440 1656.030 ;
        RECT 157.840 1472.930 159.440 1476.030 ;
        RECT 157.840 1292.930 159.440 1296.030 ;
        RECT 157.840 1112.930 159.440 1116.030 ;
        RECT 157.840 932.930 159.440 936.030 ;
        RECT 157.840 752.930 159.440 756.030 ;
        RECT 157.840 572.930 159.440 576.030 ;
        RECT 157.840 392.930 159.440 396.030 ;
        RECT 157.840 212.930 159.440 216.030 ;
        RECT 157.840 32.930 159.440 36.030 ;
        RECT 207.570 -38.270 210.670 3557.950 ;
        RECT 387.570 1774.900 390.670 3557.950 ;
        RECT 311.440 1652.930 313.040 1656.030 ;
        RECT 465.040 1652.930 466.640 1656.030 ;
        RECT 311.440 1472.930 313.040 1476.030 ;
        RECT 465.040 1472.930 466.640 1476.030 ;
        RECT 311.440 1292.930 313.040 1296.030 ;
        RECT 465.040 1292.930 466.640 1296.030 ;
        RECT 311.440 1112.930 313.040 1116.030 ;
        RECT 465.040 1112.930 466.640 1116.030 ;
        RECT 311.440 932.930 313.040 936.030 ;
        RECT 465.040 932.930 466.640 936.030 ;
        RECT 311.440 752.930 313.040 756.030 ;
        RECT 465.040 752.930 466.640 756.030 ;
        RECT 311.440 572.930 313.040 576.030 ;
        RECT 465.040 572.930 466.640 576.030 ;
        RECT 311.440 392.930 313.040 396.030 ;
        RECT 465.040 392.930 466.640 396.030 ;
        RECT 311.440 212.930 313.040 216.030 ;
        RECT 465.040 212.930 466.640 216.030 ;
        RECT 311.440 32.930 313.040 36.030 ;
        RECT 465.040 32.930 466.640 36.030 ;
        RECT 567.570 -38.270 570.670 3557.950 ;
        RECT 618.640 1652.930 620.240 1656.030 ;
        RECT 618.640 1472.930 620.240 1476.030 ;
        RECT 618.640 1292.930 620.240 1296.030 ;
        RECT 618.640 1112.930 620.240 1116.030 ;
        RECT 618.640 932.930 620.240 936.030 ;
        RECT 618.640 752.930 620.240 756.030 ;
        RECT 618.640 572.930 620.240 576.030 ;
        RECT 618.640 392.930 620.240 396.030 ;
        RECT 618.640 212.930 620.240 216.030 ;
        RECT 618.640 32.930 620.240 36.030 ;
        RECT 747.570 -38.270 750.670 3557.950 ;
        RECT 927.570 1774.900 930.670 3557.950 ;
        RECT 772.240 1652.930 773.840 1656.030 ;
        RECT 925.840 1652.930 927.440 1656.030 ;
        RECT 1079.440 1652.930 1081.040 1656.030 ;
        RECT 772.240 1472.930 773.840 1476.030 ;
        RECT 925.840 1472.930 927.440 1476.030 ;
        RECT 1079.440 1472.930 1081.040 1476.030 ;
        RECT 772.240 1292.930 773.840 1296.030 ;
        RECT 925.840 1292.930 927.440 1296.030 ;
        RECT 1079.440 1292.930 1081.040 1296.030 ;
        RECT 772.240 1112.930 773.840 1116.030 ;
        RECT 925.840 1112.930 927.440 1116.030 ;
        RECT 1079.440 1112.930 1081.040 1116.030 ;
        RECT 772.240 932.930 773.840 936.030 ;
        RECT 925.840 932.930 927.440 936.030 ;
        RECT 1079.440 932.930 1081.040 936.030 ;
        RECT 772.240 752.930 773.840 756.030 ;
        RECT 925.840 752.930 927.440 756.030 ;
        RECT 1079.440 752.930 1081.040 756.030 ;
        RECT 772.240 572.930 773.840 576.030 ;
        RECT 925.840 572.930 927.440 576.030 ;
        RECT 1079.440 572.930 1081.040 576.030 ;
        RECT 772.240 392.930 773.840 396.030 ;
        RECT 925.840 392.930 927.440 396.030 ;
        RECT 1079.440 392.930 1081.040 396.030 ;
        RECT 772.240 212.930 773.840 216.030 ;
        RECT 925.840 212.930 927.440 216.030 ;
        RECT 1079.440 212.930 1081.040 216.030 ;
        RECT 772.240 32.930 773.840 36.030 ;
        RECT 925.840 32.930 927.440 36.030 ;
        RECT 1079.440 32.930 1081.040 36.030 ;
        RECT 1107.570 -38.270 1110.670 3557.950 ;
        RECT 1233.040 1652.930 1234.640 1656.030 ;
        RECT 1233.040 1472.930 1234.640 1476.030 ;
        RECT 1233.040 1292.930 1234.640 1296.030 ;
        RECT 1233.040 1112.930 1234.640 1116.030 ;
        RECT 1233.040 932.930 1234.640 936.030 ;
        RECT 1233.040 752.930 1234.640 756.030 ;
        RECT 1233.040 572.930 1234.640 576.030 ;
        RECT 1233.040 392.930 1234.640 396.030 ;
        RECT 1233.040 212.930 1234.640 216.030 ;
        RECT 1233.040 32.930 1234.640 36.030 ;
        RECT 1287.570 -38.270 1290.670 3557.950 ;
        RECT 1386.640 1652.930 1388.240 1656.030 ;
        RECT 1386.640 1472.930 1388.240 1476.030 ;
        RECT 1386.640 1292.930 1388.240 1296.030 ;
        RECT 1386.640 1112.930 1388.240 1116.030 ;
        RECT 1386.640 932.930 1388.240 936.030 ;
        RECT 1386.640 752.930 1388.240 756.030 ;
        RECT 1386.640 572.930 1388.240 576.030 ;
        RECT 1386.640 392.930 1388.240 396.030 ;
        RECT 1386.640 212.930 1388.240 216.030 ;
        RECT 1386.640 32.930 1388.240 36.030 ;
        RECT 1467.570 -38.270 1470.670 3557.950 ;
        RECT 1540.240 1652.930 1541.840 1656.030 ;
        RECT 1540.240 1472.930 1541.840 1476.030 ;
        RECT 1540.240 1292.930 1541.840 1296.030 ;
        RECT 1540.240 1112.930 1541.840 1116.030 ;
        RECT 1540.240 932.930 1541.840 936.030 ;
        RECT 1540.240 752.930 1541.840 756.030 ;
        RECT 1540.240 572.930 1541.840 576.030 ;
        RECT 1540.240 392.930 1541.840 396.030 ;
        RECT 1540.240 212.930 1541.840 216.030 ;
        RECT 1540.240 32.930 1541.840 36.030 ;
        RECT 1647.570 -38.270 1650.670 3557.950 ;
        RECT 1693.840 1652.930 1695.440 1656.030 ;
        RECT 1693.840 1472.930 1695.440 1476.030 ;
        RECT 1693.840 1292.930 1695.440 1296.030 ;
        RECT 1693.840 1112.930 1695.440 1116.030 ;
        RECT 1693.840 932.930 1695.440 936.030 ;
        RECT 1693.840 752.930 1695.440 756.030 ;
        RECT 1693.840 572.930 1695.440 576.030 ;
        RECT 1693.840 392.930 1695.440 396.030 ;
        RECT 1693.840 212.930 1695.440 216.030 ;
        RECT 1693.840 32.930 1695.440 36.030 ;
        RECT 1827.570 -38.270 1830.670 3557.950 ;
        RECT 1847.440 1652.930 1849.040 1656.030 ;
        RECT 2001.040 1652.930 2002.640 1656.030 ;
        RECT 1847.440 1472.930 1849.040 1476.030 ;
        RECT 2001.040 1472.930 2002.640 1476.030 ;
        RECT 1847.440 1292.930 1849.040 1296.030 ;
        RECT 2001.040 1292.930 2002.640 1296.030 ;
        RECT 1847.440 1112.930 1849.040 1116.030 ;
        RECT 2001.040 1112.930 2002.640 1116.030 ;
        RECT 1847.440 932.930 1849.040 936.030 ;
        RECT 2001.040 932.930 2002.640 936.030 ;
        RECT 1847.440 752.930 1849.040 756.030 ;
        RECT 2001.040 752.930 2002.640 756.030 ;
        RECT 1847.440 572.930 1849.040 576.030 ;
        RECT 2001.040 572.930 2002.640 576.030 ;
        RECT 1847.440 392.930 1849.040 396.030 ;
        RECT 2001.040 392.930 2002.640 396.030 ;
        RECT 1847.440 212.930 1849.040 216.030 ;
        RECT 2001.040 212.930 2002.640 216.030 ;
        RECT 1847.440 32.930 1849.040 36.030 ;
        RECT 2001.040 32.930 2002.640 36.030 ;
        RECT 2007.570 -38.270 2010.670 3557.950 ;
        RECT 2154.640 1652.930 2156.240 1656.030 ;
        RECT 2154.640 1472.930 2156.240 1476.030 ;
        RECT 2154.640 1292.930 2156.240 1296.030 ;
        RECT 2154.640 1112.930 2156.240 1116.030 ;
        RECT 2154.640 932.930 2156.240 936.030 ;
        RECT 2154.640 752.930 2156.240 756.030 ;
        RECT 2154.640 572.930 2156.240 576.030 ;
        RECT 2154.640 392.930 2156.240 396.030 ;
        RECT 2154.640 212.930 2156.240 216.030 ;
        RECT 2154.640 32.930 2156.240 36.030 ;
        RECT 2187.570 -38.270 2190.670 3557.950 ;
        RECT 2308.240 1652.930 2309.840 1656.030 ;
        RECT 2308.240 1472.930 2309.840 1476.030 ;
        RECT 2308.240 1292.930 2309.840 1296.030 ;
        RECT 2308.240 1112.930 2309.840 1116.030 ;
        RECT 2308.240 932.930 2309.840 936.030 ;
        RECT 2308.240 752.930 2309.840 756.030 ;
        RECT 2308.240 572.930 2309.840 576.030 ;
        RECT 2308.240 392.930 2309.840 396.030 ;
        RECT 2308.240 212.930 2309.840 216.030 ;
        RECT 2308.240 32.930 2309.840 36.030 ;
        RECT 2367.570 -38.270 2370.670 3557.950 ;
        RECT 2461.840 1652.930 2463.440 1656.030 ;
        RECT 2461.840 1472.930 2463.440 1476.030 ;
        RECT 2461.840 1292.930 2463.440 1296.030 ;
        RECT 2461.840 1112.930 2463.440 1116.030 ;
        RECT 2461.840 932.930 2463.440 936.030 ;
        RECT 2461.840 752.930 2463.440 756.030 ;
        RECT 2461.840 572.930 2463.440 576.030 ;
        RECT 2461.840 392.930 2463.440 396.030 ;
        RECT 2461.840 212.930 2463.440 216.030 ;
        RECT 2461.840 32.930 2463.440 36.030 ;
        RECT 2547.570 -38.270 2550.670 3557.950 ;
        RECT 2615.440 1652.930 2617.040 1656.030 ;
        RECT 2615.440 1472.930 2617.040 1476.030 ;
        RECT 2615.440 1292.930 2617.040 1296.030 ;
        RECT 2615.440 1112.930 2617.040 1116.030 ;
        RECT 2615.440 932.930 2617.040 936.030 ;
        RECT 2615.440 752.930 2617.040 756.030 ;
        RECT 2615.440 572.930 2617.040 576.030 ;
        RECT 2615.440 392.930 2617.040 396.030 ;
        RECT 2615.440 212.930 2617.040 216.030 ;
        RECT 2615.440 32.930 2617.040 36.030 ;
        RECT 2727.570 -38.270 2730.670 3557.950 ;
        RECT 2769.040 1652.930 2770.640 1656.030 ;
        RECT 2769.040 1472.930 2770.640 1476.030 ;
        RECT 2769.040 1292.930 2770.640 1296.030 ;
        RECT 2769.040 1112.930 2770.640 1116.030 ;
        RECT 2769.040 932.930 2770.640 936.030 ;
        RECT 2769.040 752.930 2770.640 756.030 ;
        RECT 2769.040 572.930 2770.640 576.030 ;
        RECT 2769.040 392.930 2770.640 396.030 ;
        RECT 2769.040 212.930 2770.640 216.030 ;
        RECT 2769.040 32.930 2770.640 36.030 ;
        RECT 2907.570 -38.270 2910.670 3557.950 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -43.630 3452.930 2963.250 3456.030 ;
        RECT -43.630 3272.930 2963.250 3276.030 ;
        RECT -43.630 3092.930 2963.250 3096.030 ;
        RECT -43.630 2912.930 2963.250 2916.030 ;
        RECT -43.630 2732.930 2963.250 2736.030 ;
        RECT -43.630 2552.930 2963.250 2556.030 ;
        RECT -43.630 2372.930 2963.250 2376.030 ;
        RECT -43.630 2192.930 2963.250 2196.030 ;
        RECT -43.630 2012.930 2963.250 2016.030 ;
        RECT -43.630 1832.930 2963.250 1836.030 ;
        RECT -43.630 1652.930 2963.250 1656.030 ;
        RECT -43.630 1472.930 2963.250 1476.030 ;
        RECT -43.630 1292.930 2963.250 1296.030 ;
        RECT -43.630 1112.930 2963.250 1116.030 ;
        RECT -43.630 932.930 2963.250 936.030 ;
        RECT -43.630 752.930 2963.250 756.030 ;
        RECT -43.630 572.930 2963.250 576.030 ;
        RECT -43.630 392.930 2963.250 396.030 ;
        RECT -43.630 212.930 2963.250 216.030 ;
        RECT -43.630 32.930 2963.250 36.030 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
        RECT 244.770 -38.270 247.870 3557.950 ;
        RECT 424.770 -38.270 427.870 3557.950 ;
        RECT 604.770 -38.270 607.870 3557.950 ;
        RECT 784.770 -38.270 787.870 3557.950 ;
        RECT 964.770 -38.270 967.870 3557.950 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
        RECT -43.630 970.130 2963.250 973.230 ;
        RECT -43.630 790.130 2963.250 793.230 ;
        RECT -43.630 610.130 2963.250 613.230 ;
        RECT -43.630 430.130 2963.250 433.230 ;
        RECT -43.630 250.130 2963.250 253.230 ;
        RECT -43.630 70.130 2963.250 73.230 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.050 14.010 102.190 15.300 ;
        RECT 101.820 13.870 102.190 14.010 ;
        RECT 1.930 0.410 2.210 0.525 ;
        RECT 2.710 0.410 3.270 2.400 ;
        RECT 101.820 0.525 101.960 13.870 ;
        RECT 1.930 0.270 3.270 0.410 ;
        RECT 1.930 0.155 2.210 0.270 ;
        RECT 2.710 -4.800 3.270 0.270 ;
        RECT 101.750 0.155 102.030 0.525 ;
      LAYER met3 ;
        RECT 1.905 0.490 2.235 0.505 ;
        RECT 101.725 0.490 102.055 0.505 ;
        RECT 1.905 0.190 102.055 0.490 ;
        RECT 1.905 0.175 2.235 0.190 ;
        RECT 101.725 0.175 102.055 0.190 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.570 14.010 107.710 15.300 ;
        RECT 107.340 13.870 107.710 14.010 ;
        RECT 7.450 1.090 7.730 1.205 ;
        RECT 8.230 1.090 8.790 2.400 ;
        RECT 107.340 1.205 107.480 13.870 ;
        RECT 7.450 0.950 8.790 1.090 ;
        RECT 7.450 0.835 7.730 0.950 ;
        RECT 8.230 -4.800 8.790 0.950 ;
        RECT 107.270 0.835 107.550 1.205 ;
      LAYER met3 ;
        RECT 7.425 1.170 7.755 1.185 ;
        RECT 107.245 1.170 107.575 1.185 ;
        RECT 7.425 0.870 107.575 1.170 ;
        RECT 7.425 0.855 7.755 0.870 ;
        RECT 107.245 0.855 107.575 0.870 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.090 14.010 113.230 15.300 ;
        RECT 112.860 13.870 113.230 14.010 ;
        RECT 14.210 1.770 14.770 2.400 ;
        RECT 112.860 1.885 113.000 13.870 ;
        RECT 16.650 1.770 16.930 1.885 ;
        RECT 14.210 1.630 16.930 1.770 ;
        RECT 14.210 -4.800 14.770 1.630 ;
        RECT 16.650 1.515 16.930 1.630 ;
        RECT 112.790 1.515 113.070 1.885 ;
      LAYER met3 ;
        RECT 16.625 1.850 16.955 1.865 ;
        RECT 112.765 1.850 113.095 1.865 ;
        RECT 16.625 1.550 113.095 1.850 ;
        RECT 16.625 1.535 16.955 1.550 ;
        RECT 112.765 1.535 113.095 1.550 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.170 14.010 135.310 15.300 ;
        RECT 134.940 13.870 135.310 14.010 ;
        RECT 134.940 2.565 135.080 13.870 ;
        RECT 41.030 2.450 41.310 2.565 ;
        RECT 38.130 1.770 38.690 2.400 ;
        RECT 40.640 2.310 41.310 2.450 ;
        RECT 40.640 1.770 40.780 2.310 ;
        RECT 41.030 2.195 41.310 2.310 ;
        RECT 134.870 2.195 135.150 2.565 ;
        RECT 38.130 1.630 40.780 1.770 ;
        RECT 38.130 -4.800 38.690 1.630 ;
      LAYER met3 ;
        RECT 41.005 2.530 41.335 2.545 ;
        RECT 134.845 2.530 135.175 2.545 ;
        RECT 41.005 2.230 135.175 2.530 ;
        RECT 41.005 2.215 41.335 2.230 ;
        RECT 134.845 2.215 135.175 2.230 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 14.010 321.910 14.125 ;
        RECT 322.850 14.010 322.990 15.300 ;
        RECT 321.630 13.870 322.990 14.010 ;
        RECT 321.630 13.755 321.910 13.870 ;
        RECT 239.290 13.075 239.570 13.445 ;
        RECT 239.360 2.400 239.500 13.075 ;
        RECT 239.150 -4.800 239.710 2.400 ;
      LAYER met3 ;
        RECT 239.470 19.530 239.850 19.540 ;
        RECT 299.270 19.530 299.650 19.540 ;
        RECT 239.470 19.230 299.650 19.530 ;
        RECT 239.470 19.220 239.850 19.230 ;
        RECT 299.270 19.220 299.650 19.230 ;
        RECT 299.270 14.090 299.650 14.100 ;
        RECT 321.605 14.090 321.935 14.105 ;
        RECT 299.270 13.790 321.935 14.090 ;
        RECT 299.270 13.780 299.650 13.790 ;
        RECT 321.605 13.775 321.935 13.790 ;
        RECT 239.265 13.420 239.595 13.425 ;
        RECT 239.265 13.410 239.850 13.420 ;
        RECT 239.040 13.110 239.850 13.410 ;
        RECT 239.265 13.100 239.850 13.110 ;
        RECT 239.265 13.095 239.595 13.100 ;
      LAYER met4 ;
        RECT 239.495 19.215 239.825 19.545 ;
        RECT 299.295 19.215 299.625 19.545 ;
        RECT 239.510 13.425 239.810 19.215 ;
        RECT 299.310 14.105 299.610 19.215 ;
        RECT 299.295 13.775 299.625 14.105 ;
        RECT 239.495 13.095 239.825 13.425 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 256.750 14.180 257.070 14.240 ;
        RECT 296.310 14.180 296.630 14.240 ;
        RECT 256.750 14.040 296.630 14.180 ;
        RECT 256.750 13.980 257.070 14.040 ;
        RECT 296.310 13.980 296.630 14.040 ;
        RECT 296.310 6.700 296.630 6.760 ;
        RECT 339.090 6.700 339.410 6.760 ;
        RECT 296.310 6.560 339.410 6.700 ;
        RECT 296.310 6.500 296.630 6.560 ;
        RECT 339.090 6.500 339.410 6.560 ;
      LAYER met2 ;
        RECT 256.780 13.950 257.040 14.270 ;
        RECT 296.340 13.950 296.600 14.270 ;
        RECT 339.410 14.010 339.550 15.300 ;
        RECT 256.840 2.400 256.980 13.950 ;
        RECT 296.400 6.790 296.540 13.950 ;
        RECT 339.180 13.870 339.550 14.010 ;
        RECT 339.180 6.790 339.320 13.870 ;
        RECT 296.340 6.470 296.600 6.790 ;
        RECT 339.120 6.470 339.380 6.790 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 275.610 0.920 275.930 0.980 ;
        RECT 355.650 0.920 355.970 0.980 ;
        RECT 275.610 0.780 355.970 0.920 ;
        RECT 275.610 0.720 275.930 0.780 ;
        RECT 355.650 0.720 355.970 0.780 ;
      LAYER met2 ;
        RECT 355.970 14.010 356.110 15.300 ;
        RECT 355.740 13.870 356.110 14.010 ;
        RECT 274.570 1.090 275.130 2.400 ;
        RECT 274.570 1.010 275.840 1.090 ;
        RECT 355.740 1.010 355.880 13.870 ;
        RECT 274.570 0.950 275.900 1.010 ;
        RECT 274.570 -4.800 275.130 0.950 ;
        RECT 275.640 0.690 275.900 0.950 ;
        RECT 355.680 0.690 355.940 1.010 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.530 14.805 372.670 15.300 ;
        RECT 372.460 14.435 372.740 14.805 ;
        RECT 292.190 13.755 292.470 14.125 ;
        RECT 292.260 2.400 292.400 13.755 ;
        RECT 292.050 -4.800 292.610 2.400 ;
      LAYER met3 ;
        RECT 292.870 14.470 324.450 14.770 ;
        RECT 292.165 14.090 292.495 14.105 ;
        RECT 292.870 14.090 293.170 14.470 ;
        RECT 292.165 13.790 293.170 14.090 ;
        RECT 324.150 14.090 324.450 14.470 ;
        RECT 372.435 14.455 372.765 14.785 ;
        RECT 372.450 14.090 372.750 14.455 ;
        RECT 324.150 13.790 372.750 14.090 ;
        RECT 292.165 13.775 292.495 13.790 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 309.190 2.280 309.510 2.340 ;
        RECT 388.770 2.280 389.090 2.340 ;
        RECT 309.190 2.140 389.090 2.280 ;
        RECT 309.190 2.080 309.510 2.140 ;
        RECT 388.770 2.080 389.090 2.140 ;
      LAYER met2 ;
        RECT 389.090 14.010 389.230 15.300 ;
        RECT 388.860 13.870 389.230 14.010 ;
        RECT 309.220 2.050 309.480 2.370 ;
        RECT 309.280 1.770 309.420 2.050 ;
        RECT 309.990 1.770 310.550 2.400 ;
        RECT 388.860 2.370 389.000 13.870 ;
        RECT 388.800 2.050 389.060 2.370 ;
        RECT 309.280 1.630 310.550 1.770 ;
        RECT 309.990 -4.800 310.550 1.630 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.650 14.010 405.790 15.300 ;
        RECT 405.420 13.870 405.790 14.010 ;
        RECT 405.420 10.725 405.560 13.870 ;
        RECT 327.610 10.355 327.890 10.725 ;
        RECT 405.350 10.355 405.630 10.725 ;
        RECT 327.680 2.400 327.820 10.355 ;
        RECT 327.470 -4.800 328.030 2.400 ;
      LAYER met3 ;
        RECT 327.585 10.690 327.915 10.705 ;
        RECT 405.325 10.690 405.655 10.705 ;
        RECT 327.585 10.390 405.655 10.690 ;
        RECT 327.585 10.375 327.915 10.390 ;
        RECT 405.325 10.375 405.655 10.390 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.210 14.010 422.350 15.300 ;
        RECT 421.980 13.870 422.350 14.010 ;
        RECT 421.980 12.085 422.120 13.870 ;
        RECT 345.550 11.715 345.830 12.085 ;
        RECT 421.910 11.715 422.190 12.085 ;
        RECT 345.620 2.400 345.760 11.715 ;
        RECT 345.410 -4.800 345.970 2.400 ;
      LAYER met3 ;
        RECT 345.525 12.050 345.855 12.065 ;
        RECT 421.885 12.050 422.215 12.065 ;
        RECT 345.525 11.750 422.215 12.050 ;
        RECT 345.525 11.735 345.855 11.750 ;
        RECT 421.885 11.735 422.215 11.750 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.770 14.010 438.910 15.300 ;
        RECT 438.540 13.870 438.910 14.010 ;
        RECT 438.540 12.765 438.680 13.870 ;
        RECT 363.030 12.395 363.310 12.765 ;
        RECT 438.470 12.395 438.750 12.765 ;
        RECT 363.100 2.400 363.240 12.395 ;
        RECT 362.890 -4.800 363.450 2.400 ;
      LAYER met3 ;
        RECT 363.005 12.730 363.335 12.745 ;
        RECT 438.445 12.730 438.775 12.745 ;
        RECT 363.005 12.430 438.775 12.730 ;
        RECT 363.005 12.415 363.335 12.430 ;
        RECT 438.445 12.415 438.775 12.430 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.330 14.125 455.470 15.300 ;
        RECT 380.970 13.755 381.250 14.125 ;
        RECT 455.260 13.755 455.540 14.125 ;
        RECT 381.040 2.400 381.180 13.755 ;
        RECT 380.830 -4.800 381.390 2.400 ;
      LAYER met3 ;
        RECT 380.945 14.090 381.275 14.105 ;
        RECT 455.235 14.090 455.565 14.105 ;
        RECT 380.945 13.790 455.565 14.090 ;
        RECT 380.945 13.775 381.275 13.790 ;
        RECT 455.235 13.775 455.565 13.790 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 397.510 1.600 397.830 1.660 ;
        RECT 471.570 1.600 471.890 1.660 ;
        RECT 397.510 1.460 471.890 1.600 ;
        RECT 397.510 1.400 397.830 1.460 ;
        RECT 471.570 1.400 471.890 1.460 ;
      LAYER met2 ;
        RECT 471.890 14.010 472.030 15.300 ;
        RECT 471.660 13.870 472.030 14.010 ;
        RECT 398.310 1.770 398.870 2.400 ;
        RECT 397.600 1.690 398.870 1.770 ;
        RECT 471.660 1.690 471.800 13.870 ;
        RECT 397.540 1.630 398.870 1.690 ;
        RECT 397.540 1.370 397.800 1.630 ;
        RECT 398.310 -4.800 398.870 1.630 ;
        RECT 471.600 1.370 471.860 1.690 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 96.210 5.340 96.530 5.400 ;
        RECT 156.930 5.340 157.250 5.400 ;
        RECT 96.210 5.200 157.250 5.340 ;
        RECT 96.210 5.140 96.530 5.200 ;
        RECT 156.930 5.140 157.250 5.200 ;
      LAYER met2 ;
        RECT 157.250 14.010 157.390 15.300 ;
        RECT 157.020 13.870 157.390 14.010 ;
        RECT 157.020 5.430 157.160 13.870 ;
        RECT 96.240 5.285 96.500 5.430 ;
        RECT 61.730 4.915 62.010 5.285 ;
        RECT 96.230 4.915 96.510 5.285 ;
        RECT 156.960 5.110 157.220 5.430 ;
        RECT 61.800 2.400 61.940 4.915 ;
        RECT 61.590 -4.800 62.150 2.400 ;
      LAYER met3 ;
        RECT 61.705 5.250 62.035 5.265 ;
        RECT 96.205 5.250 96.535 5.265 ;
        RECT 61.705 4.950 96.535 5.250 ;
        RECT 61.705 4.935 62.035 4.950 ;
        RECT 96.205 4.935 96.535 4.950 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.450 14.010 488.590 15.300 ;
        RECT 488.220 13.870 488.590 14.010 ;
        RECT 416.460 2.990 417.520 3.130 ;
        RECT 416.460 2.400 416.600 2.990 ;
        RECT 417.380 2.565 417.520 2.990 ;
        RECT 488.220 2.565 488.360 13.870 ;
        RECT 416.250 -4.800 416.810 2.400 ;
        RECT 417.310 2.195 417.590 2.565 ;
        RECT 488.150 2.195 488.430 2.565 ;
      LAYER met3 ;
        RECT 417.285 2.530 417.615 2.545 ;
        RECT 488.125 2.530 488.455 2.545 ;
        RECT 417.285 2.230 488.455 2.530 ;
        RECT 417.285 2.215 417.615 2.230 ;
        RECT 488.125 2.215 488.455 2.230 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 433.390 0.580 433.710 0.640 ;
        RECT 504.230 0.580 504.550 0.640 ;
        RECT 433.390 0.440 504.550 0.580 ;
        RECT 433.390 0.380 433.710 0.440 ;
        RECT 504.230 0.380 504.550 0.440 ;
      LAYER met2 ;
        RECT 505.010 14.010 505.150 15.300 ;
        RECT 504.320 13.870 505.150 14.010 ;
        RECT 433.420 0.410 433.680 0.670 ;
        RECT 434.190 0.410 434.750 2.400 ;
        RECT 504.320 0.670 504.460 13.870 ;
        RECT 433.420 0.350 434.750 0.410 ;
        RECT 504.260 0.350 504.520 0.670 ;
        RECT 433.480 0.270 434.750 0.350 ;
        RECT 434.190 -4.800 434.750 0.270 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.570 14.010 521.710 15.300 ;
        RECT 520.880 13.870 521.710 14.010 ;
        RECT 450.890 0.410 451.170 0.525 ;
        RECT 451.670 0.410 452.230 2.400 ;
        RECT 520.880 0.525 521.020 13.870 ;
        RECT 450.890 0.270 452.230 0.410 ;
        RECT 450.890 0.155 451.170 0.270 ;
        RECT 451.670 -4.800 452.230 0.270 ;
        RECT 520.810 0.155 521.090 0.525 ;
      LAYER met3 ;
        RECT 450.865 0.490 451.195 0.505 ;
        RECT 520.785 0.490 521.115 0.505 ;
        RECT 450.865 0.190 521.115 0.490 ;
        RECT 450.865 0.175 451.195 0.190 ;
        RECT 520.785 0.175 521.115 0.190 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.130 14.010 538.270 15.300 ;
        RECT 537.900 13.870 538.270 14.010 ;
        RECT 537.900 10.045 538.040 13.870 ;
        RECT 469.750 9.675 470.030 10.045 ;
        RECT 537.830 9.675 538.110 10.045 ;
        RECT 469.820 2.400 469.960 9.675 ;
        RECT 469.610 -4.800 470.170 2.400 ;
      LAYER met3 ;
        RECT 469.725 10.010 470.055 10.025 ;
        RECT 537.805 10.010 538.135 10.025 ;
        RECT 469.725 9.710 538.135 10.010 ;
        RECT 469.725 9.695 470.055 9.710 ;
        RECT 537.805 9.695 538.135 9.710 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.510 6.020 489.830 6.080 ;
        RECT 554.370 6.020 554.690 6.080 ;
        RECT 489.510 5.880 554.690 6.020 ;
        RECT 489.510 5.820 489.830 5.880 ;
        RECT 554.370 5.820 554.690 5.880 ;
      LAYER met2 ;
        RECT 554.690 14.010 554.830 15.300 ;
        RECT 554.460 13.870 554.830 14.010 ;
        RECT 554.460 6.110 554.600 13.870 ;
        RECT 489.540 5.790 489.800 6.110 ;
        RECT 554.400 5.790 554.660 6.110 ;
        RECT 487.090 1.770 487.650 2.400 ;
        RECT 489.600 1.770 489.740 5.790 ;
        RECT 487.090 1.630 489.740 1.770 ;
        RECT 487.090 -4.800 487.650 1.630 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.250 14.010 571.390 15.300 ;
        RECT 571.020 13.870 571.390 14.010 ;
        RECT 571.020 10.725 571.160 13.870 ;
        RECT 505.170 10.355 505.450 10.725 ;
        RECT 570.950 10.355 571.230 10.725 ;
        RECT 505.240 2.400 505.380 10.355 ;
        RECT 505.030 -4.800 505.590 2.400 ;
      LAYER met3 ;
        RECT 505.145 10.690 505.475 10.705 ;
        RECT 570.925 10.690 571.255 10.705 ;
        RECT 505.145 10.390 571.255 10.690 ;
        RECT 505.145 10.375 505.475 10.390 ;
        RECT 570.925 10.375 571.255 10.390 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.630 6.700 522.950 6.760 ;
        RECT 587.490 6.700 587.810 6.760 ;
        RECT 522.630 6.560 587.810 6.700 ;
        RECT 522.630 6.500 522.950 6.560 ;
        RECT 587.490 6.500 587.810 6.560 ;
      LAYER met2 ;
        RECT 587.810 14.010 587.950 15.300 ;
        RECT 587.580 13.870 587.950 14.010 ;
        RECT 587.580 6.790 587.720 13.870 ;
        RECT 522.660 6.470 522.920 6.790 ;
        RECT 587.520 6.470 587.780 6.790 ;
        RECT 522.720 2.400 522.860 6.470 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.370 14.010 604.510 15.300 ;
        RECT 604.140 13.870 604.510 14.010 ;
        RECT 604.140 10.045 604.280 13.870 ;
        RECT 540.590 9.675 540.870 10.045 ;
        RECT 604.070 9.675 604.350 10.045 ;
        RECT 540.660 2.400 540.800 9.675 ;
        RECT 540.450 -4.800 541.010 2.400 ;
      LAYER met3 ;
        RECT 540.565 10.010 540.895 10.025 ;
        RECT 604.045 10.010 604.375 10.025 ;
        RECT 540.565 9.710 604.375 10.010 ;
        RECT 540.565 9.695 540.895 9.710 ;
        RECT 604.045 9.695 604.375 9.710 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.930 14.010 621.070 15.300 ;
        RECT 620.700 13.870 621.070 14.010 ;
        RECT 620.700 9.365 620.840 13.870 ;
        RECT 558.070 8.995 558.350 9.365 ;
        RECT 620.630 8.995 620.910 9.365 ;
        RECT 558.140 2.400 558.280 8.995 ;
        RECT 557.930 -4.800 558.490 2.400 ;
      LAYER met3 ;
        RECT 558.045 9.330 558.375 9.345 ;
        RECT 620.605 9.330 620.935 9.345 ;
        RECT 558.045 9.030 620.935 9.330 ;
        RECT 558.045 9.015 558.375 9.030 ;
        RECT 620.605 9.015 620.935 9.030 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.490 14.010 637.630 15.300 ;
        RECT 637.260 13.870 637.630 14.010 ;
        RECT 637.260 10.725 637.400 13.870 ;
        RECT 576.010 10.355 576.290 10.725 ;
        RECT 637.190 10.355 637.470 10.725 ;
        RECT 576.080 2.400 576.220 10.355 ;
        RECT 575.870 -4.800 576.430 2.400 ;
      LAYER met3 ;
        RECT 575.985 10.690 576.315 10.705 ;
        RECT 637.165 10.690 637.495 10.705 ;
        RECT 575.985 10.390 637.495 10.690 ;
        RECT 575.985 10.375 576.315 10.390 ;
        RECT 637.165 10.375 637.495 10.390 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.330 14.805 179.470 15.300 ;
        RECT 179.260 14.435 179.540 14.805 ;
        RECT 85.190 13.755 85.470 14.125 ;
        RECT 85.260 2.400 85.400 13.755 ;
        RECT 85.050 -4.800 85.610 2.400 ;
      LAYER met3 ;
        RECT 179.235 14.770 179.565 14.785 ;
        RECT 85.870 14.470 179.565 14.770 ;
        RECT 85.165 14.090 85.495 14.105 ;
        RECT 85.870 14.090 86.170 14.470 ;
        RECT 179.235 14.455 179.565 14.470 ;
        RECT 85.165 13.790 86.170 14.090 ;
        RECT 85.165 13.775 85.495 13.790 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.050 14.010 654.190 15.300 ;
        RECT 653.820 13.870 654.190 14.010 ;
        RECT 653.820 2.565 653.960 13.870 ;
        RECT 593.810 0.410 594.370 2.400 ;
        RECT 653.750 2.195 654.030 2.565 ;
        RECT 595.790 0.410 596.070 0.525 ;
        RECT 593.810 0.270 596.070 0.410 ;
        RECT 593.810 -4.800 594.370 0.270 ;
        RECT 595.790 0.155 596.070 0.270 ;
      LAYER met3 ;
        RECT 653.725 2.530 654.055 2.545 ;
        RECT 613.950 2.230 654.055 2.530 ;
        RECT 595.765 0.490 596.095 0.505 ;
        RECT 613.950 0.490 614.250 2.230 ;
        RECT 653.725 2.215 654.055 2.230 ;
        RECT 595.765 0.190 614.250 0.490 ;
        RECT 595.765 0.175 596.095 0.190 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 612.790 0.580 613.110 0.640 ;
        RECT 669.830 0.580 670.150 0.640 ;
        RECT 612.790 0.440 670.150 0.580 ;
        RECT 612.790 0.380 613.110 0.440 ;
        RECT 669.830 0.380 670.150 0.440 ;
      LAYER met2 ;
        RECT 670.610 14.010 670.750 15.300 ;
        RECT 669.920 13.870 670.750 14.010 ;
        RECT 611.290 0.410 611.850 2.400 ;
        RECT 669.920 0.670 670.060 13.870 ;
        RECT 612.820 0.410 613.080 0.670 ;
        RECT 611.290 0.350 613.080 0.410 ;
        RECT 669.860 0.350 670.120 0.670 ;
        RECT 611.290 0.270 613.020 0.350 ;
        RECT 611.290 -4.800 611.850 0.270 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 119.210 6.020 119.530 6.080 ;
        RECT 201.090 6.020 201.410 6.080 ;
        RECT 119.210 5.880 201.410 6.020 ;
        RECT 119.210 5.820 119.530 5.880 ;
        RECT 201.090 5.820 201.410 5.880 ;
      LAYER met2 ;
        RECT 201.410 14.010 201.550 15.300 ;
        RECT 201.180 13.870 201.550 14.010 ;
        RECT 201.180 6.110 201.320 13.870 ;
        RECT 119.240 5.790 119.500 6.110 ;
        RECT 201.120 5.790 201.380 6.110 ;
        RECT 119.300 5.285 119.440 5.790 ;
        RECT 109.110 4.915 109.390 5.285 ;
        RECT 119.230 4.915 119.510 5.285 ;
        RECT 109.180 2.400 109.320 4.915 ;
        RECT 108.970 -4.800 109.530 2.400 ;
      LAYER met3 ;
        RECT 109.085 5.250 109.415 5.265 ;
        RECT 119.205 5.250 119.535 5.265 ;
        RECT 109.085 4.950 119.535 5.250 ;
        RECT 109.085 4.935 109.415 4.950 ;
        RECT 119.205 4.935 119.535 4.950 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.490 14.010 223.630 15.300 ;
        RECT 223.260 13.870 223.630 14.010 ;
        RECT 131.650 1.090 131.930 1.205 ;
        RECT 132.430 1.090 132.990 2.400 ;
        RECT 223.260 1.205 223.400 13.870 ;
        RECT 131.650 0.950 132.990 1.090 ;
        RECT 131.650 0.835 131.930 0.950 ;
        RECT 132.430 -4.800 132.990 0.950 ;
        RECT 223.190 0.835 223.470 1.205 ;
      LAYER met3 ;
        RECT 131.625 1.170 131.955 1.185 ;
        RECT 223.165 1.170 223.495 1.185 ;
        RECT 131.625 0.870 223.495 1.170 ;
        RECT 131.625 0.855 131.955 0.870 ;
        RECT 223.165 0.855 223.495 0.870 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 150.490 14.180 150.810 14.240 ;
        RECT 185.910 14.180 186.230 14.240 ;
        RECT 150.490 14.040 186.230 14.180 ;
        RECT 150.490 13.980 150.810 14.040 ;
        RECT 185.910 13.980 186.230 14.040 ;
        RECT 185.910 6.360 186.230 6.420 ;
        RECT 239.730 6.360 240.050 6.420 ;
        RECT 185.910 6.220 240.050 6.360 ;
        RECT 185.910 6.160 186.230 6.220 ;
        RECT 239.730 6.160 240.050 6.220 ;
      LAYER met2 ;
        RECT 150.520 13.950 150.780 14.270 ;
        RECT 185.940 13.950 186.200 14.270 ;
        RECT 240.050 14.010 240.190 15.300 ;
        RECT 150.580 2.400 150.720 13.950 ;
        RECT 186.000 6.450 186.140 13.950 ;
        RECT 239.820 13.870 240.190 14.010 ;
        RECT 239.820 6.450 239.960 13.870 ;
        RECT 185.940 6.130 186.200 6.450 ;
        RECT 239.760 6.130 240.020 6.450 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 168.890 0.580 169.210 0.640 ;
        RECT 255.830 0.580 256.150 0.640 ;
        RECT 168.890 0.440 256.150 0.580 ;
        RECT 168.890 0.380 169.210 0.440 ;
        RECT 255.830 0.380 256.150 0.440 ;
      LAYER met2 ;
        RECT 256.610 14.690 256.750 15.300 ;
        RECT 255.920 14.550 256.750 14.690 ;
        RECT 168.060 2.990 169.120 3.130 ;
        RECT 168.060 2.400 168.200 2.990 ;
        RECT 167.850 -4.800 168.410 2.400 ;
        RECT 168.980 0.670 169.120 2.990 ;
        RECT 255.920 0.670 256.060 14.550 ;
        RECT 168.920 0.350 169.180 0.670 ;
        RECT 255.860 0.350 256.120 0.670 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 184.990 0.920 185.310 0.980 ;
        RECT 272.850 0.920 273.170 0.980 ;
        RECT 184.990 0.780 273.170 0.920 ;
        RECT 184.990 0.720 185.310 0.780 ;
        RECT 272.850 0.720 273.170 0.780 ;
      LAYER met2 ;
        RECT 273.170 14.010 273.310 15.300 ;
        RECT 272.940 13.870 273.310 14.010 ;
        RECT 185.790 1.090 186.350 2.400 ;
        RECT 185.080 1.010 186.350 1.090 ;
        RECT 272.940 1.010 273.080 13.870 ;
        RECT 185.020 0.950 186.350 1.010 ;
        RECT 185.020 0.690 185.280 0.950 ;
        RECT 185.790 -4.800 186.350 0.950 ;
        RECT 272.880 0.690 273.140 1.010 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.730 14.125 289.870 15.300 ;
        RECT 289.660 13.755 289.940 14.125 ;
        RECT 203.870 13.330 204.150 13.445 ;
        RECT 203.480 13.190 204.150 13.330 ;
        RECT 203.480 2.400 203.620 13.190 ;
        RECT 203.870 13.075 204.150 13.190 ;
        RECT 203.270 -4.800 203.830 2.400 ;
      LAYER met3 ;
        RECT 289.635 14.090 289.965 14.105 ;
        RECT 208.230 13.790 264.650 14.090 ;
        RECT 203.845 13.410 204.175 13.425 ;
        RECT 208.230 13.410 208.530 13.790 ;
        RECT 203.845 13.110 208.530 13.410 ;
        RECT 203.845 13.095 204.175 13.110 ;
        RECT 264.350 12.730 264.650 13.790 ;
        RECT 266.190 13.790 289.965 14.090 ;
        RECT 266.190 12.730 266.490 13.790 ;
        RECT 289.635 13.775 289.965 13.790 ;
        RECT 264.350 12.430 266.490 12.730 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.290 14.010 306.430 15.300 ;
        RECT 306.060 13.870 306.430 14.010 ;
        RECT 221.210 0.410 221.770 2.400 ;
        RECT 306.060 0.525 306.200 13.870 ;
        RECT 223.190 0.410 223.470 0.525 ;
        RECT 221.210 0.270 223.470 0.410 ;
        RECT 221.210 -4.800 221.770 0.270 ;
        RECT 223.190 0.155 223.470 0.270 ;
        RECT 305.990 0.155 306.270 0.525 ;
      LAYER met3 ;
        RECT 223.165 0.490 223.495 0.505 ;
        RECT 305.965 0.490 306.295 0.505 ;
        RECT 223.165 0.190 306.295 0.490 ;
        RECT 223.165 0.175 223.495 0.190 ;
        RECT 305.965 0.175 306.295 0.190 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 47.910 6.020 48.230 6.080 ;
        RECT 118.290 6.020 118.610 6.080 ;
        RECT 47.910 5.880 118.610 6.020 ;
        RECT 47.910 5.820 48.230 5.880 ;
        RECT 118.290 5.820 118.610 5.880 ;
      LAYER met2 ;
        RECT 118.610 14.010 118.750 15.300 ;
        RECT 118.380 13.870 118.750 14.010 ;
        RECT 118.380 6.110 118.520 13.870 ;
        RECT 47.940 5.790 48.200 6.110 ;
        RECT 118.320 5.790 118.580 6.110 ;
        RECT 48.000 3.245 48.140 5.790 ;
        RECT 20.330 2.875 20.610 3.245 ;
        RECT 47.930 2.875 48.210 3.245 ;
        RECT 20.400 2.400 20.540 2.875 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER met3 ;
        RECT 20.305 3.210 20.635 3.225 ;
        RECT 47.905 3.210 48.235 3.225 ;
        RECT 20.305 2.910 48.235 3.210 ;
        RECT 20.305 2.895 20.635 2.910 ;
        RECT 47.905 2.895 48.235 2.910 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 89.310 5.000 89.630 5.060 ;
        RECT 140.370 5.000 140.690 5.060 ;
        RECT 89.310 4.860 140.690 5.000 ;
        RECT 89.310 4.800 89.630 4.860 ;
        RECT 140.370 4.800 140.690 4.860 ;
      LAYER met2 ;
        RECT 140.690 14.010 140.830 15.300 ;
        RECT 140.460 13.870 140.830 14.010 ;
        RECT 140.460 5.090 140.600 13.870 ;
        RECT 89.340 4.770 89.600 5.090 ;
        RECT 140.400 4.770 140.660 5.090 ;
        RECT 89.400 3.925 89.540 4.770 ;
        RECT 43.790 3.555 44.070 3.925 ;
        RECT 89.330 3.555 89.610 3.925 ;
        RECT 43.860 2.400 44.000 3.555 ;
        RECT 43.650 -4.800 44.210 2.400 ;
      LAYER met3 ;
        RECT 43.765 3.890 44.095 3.905 ;
        RECT 89.305 3.890 89.635 3.905 ;
        RECT 43.765 3.590 89.635 3.890 ;
        RECT 43.765 3.575 44.095 3.590 ;
        RECT 89.305 3.575 89.635 3.590 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 243.870 1.940 244.190 2.000 ;
        RECT 328.510 1.940 328.830 2.000 ;
        RECT 243.870 1.800 328.830 1.940 ;
        RECT 243.870 1.740 244.190 1.800 ;
        RECT 328.510 1.740 328.830 1.800 ;
      LAYER met2 ;
        RECT 328.370 14.010 328.510 15.300 ;
        RECT 328.370 13.870 328.740 14.010 ;
        RECT 243.900 1.770 244.160 2.030 ;
        RECT 244.670 1.770 245.230 2.400 ;
        RECT 328.600 2.030 328.740 13.870 ;
        RECT 243.900 1.710 245.230 1.770 ;
        RECT 328.540 1.710 328.800 2.030 ;
        RECT 243.960 1.630 245.230 1.710 ;
        RECT 244.670 -4.800 245.230 1.630 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.930 14.805 345.070 15.300 ;
        RECT 344.860 14.435 345.140 14.805 ;
        RECT 265.050 13.075 265.330 13.445 ;
        RECT 262.610 1.770 263.170 2.400 ;
        RECT 265.120 1.770 265.260 13.075 ;
        RECT 262.610 1.630 265.260 1.770 ;
        RECT 262.610 -4.800 263.170 1.630 ;
      LAYER met3 ;
        RECT 275.850 15.150 334.570 15.450 ;
        RECT 275.850 14.770 276.150 15.150 ;
        RECT 265.270 14.470 276.150 14.770 ;
        RECT 334.270 14.770 334.570 15.150 ;
        RECT 344.835 14.770 345.165 14.785 ;
        RECT 334.270 14.470 345.165 14.770 ;
        RECT 265.270 13.425 265.570 14.470 ;
        RECT 344.835 14.455 345.165 14.470 ;
        RECT 265.025 13.110 265.570 13.425 ;
        RECT 265.025 13.095 265.355 13.110 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.050 1.260 282.370 1.320 ;
        RECT 361.170 1.260 361.490 1.320 ;
        RECT 282.050 1.120 361.490 1.260 ;
        RECT 282.050 1.060 282.370 1.120 ;
        RECT 361.170 1.060 361.490 1.120 ;
      LAYER met2 ;
        RECT 361.490 14.010 361.630 15.300 ;
        RECT 361.260 13.870 361.630 14.010 ;
        RECT 280.090 1.090 280.650 2.400 ;
        RECT 361.260 1.350 361.400 13.870 ;
        RECT 282.080 1.090 282.340 1.350 ;
        RECT 280.090 1.030 282.340 1.090 ;
        RECT 361.200 1.030 361.460 1.350 ;
        RECT 280.090 0.950 282.280 1.030 ;
        RECT 280.090 -4.800 280.650 0.950 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.050 14.010 378.190 15.300 ;
        RECT 377.820 13.870 378.190 14.010 ;
        RECT 377.820 10.045 377.960 13.870 ;
        RECT 298.170 9.675 298.450 10.045 ;
        RECT 377.750 9.675 378.030 10.045 ;
        RECT 298.240 2.400 298.380 9.675 ;
        RECT 298.030 -4.800 298.590 2.400 ;
      LAYER met3 ;
        RECT 298.145 10.010 298.475 10.025 ;
        RECT 377.725 10.010 378.055 10.025 ;
        RECT 298.145 9.710 378.055 10.010 ;
        RECT 298.145 9.695 298.475 9.710 ;
        RECT 377.725 9.695 378.055 9.710 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.010 2.620 317.330 2.680 ;
        RECT 394.290 2.620 394.610 2.680 ;
        RECT 317.010 2.480 394.610 2.620 ;
        RECT 317.010 2.420 317.330 2.480 ;
        RECT 394.290 2.420 394.610 2.480 ;
      LAYER met2 ;
        RECT 394.610 14.010 394.750 15.300 ;
        RECT 394.380 13.870 394.750 14.010 ;
        RECT 394.380 2.710 394.520 13.870 ;
        RECT 315.970 1.770 316.530 2.400 ;
        RECT 317.040 2.390 317.300 2.710 ;
        RECT 394.320 2.390 394.580 2.710 ;
        RECT 317.100 1.770 317.240 2.390 ;
        RECT 315.970 1.630 317.240 1.770 ;
        RECT 315.970 -4.800 316.530 1.630 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.170 14.010 411.310 15.300 ;
        RECT 410.940 13.870 411.310 14.010 ;
        RECT 410.940 11.405 411.080 13.870 ;
        RECT 334.970 11.290 335.250 11.405 ;
        RECT 334.120 11.150 335.250 11.290 ;
        RECT 334.120 3.130 334.260 11.150 ;
        RECT 334.970 11.035 335.250 11.150 ;
        RECT 410.870 11.035 411.150 11.405 ;
        RECT 333.660 2.990 334.260 3.130 ;
        RECT 333.660 2.400 333.800 2.990 ;
        RECT 333.450 -4.800 334.010 2.400 ;
      LAYER met3 ;
        RECT 334.945 11.370 335.275 11.385 ;
        RECT 410.845 11.370 411.175 11.385 ;
        RECT 334.945 11.070 411.175 11.370 ;
        RECT 334.945 11.055 335.275 11.070 ;
        RECT 410.845 11.055 411.175 11.070 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.510 14.180 351.830 14.240 ;
        RECT 386.010 14.180 386.330 14.240 ;
        RECT 351.510 14.040 386.330 14.180 ;
        RECT 351.510 13.980 351.830 14.040 ;
        RECT 386.010 13.980 386.330 14.040 ;
        RECT 386.010 6.360 386.330 6.420 ;
        RECT 427.410 6.360 427.730 6.420 ;
        RECT 386.010 6.220 427.730 6.360 ;
        RECT 386.010 6.160 386.330 6.220 ;
        RECT 427.410 6.160 427.730 6.220 ;
      LAYER met2 ;
        RECT 351.540 13.950 351.800 14.270 ;
        RECT 386.040 13.950 386.300 14.270 ;
        RECT 427.730 14.010 427.870 15.300 ;
        RECT 351.600 2.400 351.740 13.950 ;
        RECT 386.100 6.450 386.240 13.950 ;
        RECT 427.500 13.870 427.870 14.010 ;
        RECT 427.500 6.450 427.640 13.870 ;
        RECT 386.040 6.130 386.300 6.450 ;
        RECT 427.440 6.130 427.700 6.450 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 368.070 0.920 368.390 0.980 ;
        RECT 443.970 0.920 444.290 0.980 ;
        RECT 368.070 0.780 444.290 0.920 ;
        RECT 368.070 0.720 368.390 0.780 ;
        RECT 443.970 0.720 444.290 0.780 ;
      LAYER met2 ;
        RECT 444.290 14.010 444.430 15.300 ;
        RECT 444.060 13.870 444.430 14.010 ;
        RECT 368.870 1.090 369.430 2.400 ;
        RECT 368.160 1.010 369.430 1.090 ;
        RECT 444.060 1.010 444.200 13.870 ;
        RECT 368.100 0.950 369.430 1.010 ;
        RECT 368.100 0.690 368.360 0.950 ;
        RECT 368.870 -4.800 369.430 0.950 ;
        RECT 444.000 0.690 444.260 1.010 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.850 14.010 460.990 15.300 ;
        RECT 460.620 13.870 460.990 14.010 ;
        RECT 460.620 3.245 460.760 13.870 ;
        RECT 386.950 2.875 387.230 3.245 ;
        RECT 460.550 2.875 460.830 3.245 ;
        RECT 387.020 2.400 387.160 2.875 ;
        RECT 386.810 -4.800 387.370 2.400 ;
      LAYER met3 ;
        RECT 386.925 3.210 387.255 3.225 ;
        RECT 460.525 3.210 460.855 3.225 ;
        RECT 386.925 2.910 460.855 3.210 ;
        RECT 386.925 2.895 387.255 2.910 ;
        RECT 460.525 2.895 460.855 2.910 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 6.020 407.490 6.080 ;
        RECT 477.090 6.020 477.410 6.080 ;
        RECT 407.170 5.880 477.410 6.020 ;
        RECT 407.170 5.820 407.490 5.880 ;
        RECT 477.090 5.820 477.410 5.880 ;
      LAYER met2 ;
        RECT 477.410 14.010 477.550 15.300 ;
        RECT 477.180 13.870 477.550 14.010 ;
        RECT 477.180 6.110 477.320 13.870 ;
        RECT 407.200 5.790 407.460 6.110 ;
        RECT 477.120 5.790 477.380 6.110 ;
        RECT 404.290 1.770 404.850 2.400 ;
        RECT 407.260 1.770 407.400 5.790 ;
        RECT 404.290 1.630 407.400 1.770 ;
        RECT 404.290 -4.800 404.850 1.630 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 68.610 0.580 68.930 0.640 ;
        RECT 162.910 0.580 163.230 0.640 ;
        RECT 68.610 0.440 163.230 0.580 ;
        RECT 68.610 0.380 68.930 0.440 ;
        RECT 162.910 0.380 163.230 0.440 ;
      LAYER met2 ;
        RECT 162.770 14.010 162.910 15.300 ;
        RECT 162.770 13.870 163.140 14.010 ;
        RECT 67.570 0.410 68.130 2.400 ;
        RECT 163.000 0.670 163.140 13.870 ;
        RECT 68.640 0.410 68.900 0.670 ;
        RECT 67.570 0.350 68.900 0.410 ;
        RECT 162.940 0.350 163.200 0.670 ;
        RECT 67.570 0.270 68.840 0.350 ;
        RECT 67.570 -4.800 68.130 0.270 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.970 14.010 494.110 15.300 ;
        RECT 493.970 13.870 494.340 14.010 ;
        RECT 422.440 2.990 423.500 3.130 ;
        RECT 422.440 2.400 422.580 2.990 ;
        RECT 422.230 -4.800 422.790 2.400 ;
        RECT 423.360 1.885 423.500 2.990 ;
        RECT 494.200 2.565 494.340 13.870 ;
        RECT 494.130 2.195 494.410 2.565 ;
        RECT 423.290 1.515 423.570 1.885 ;
      LAYER met3 ;
        RECT 494.105 2.530 494.435 2.545 ;
        RECT 494.105 2.215 494.650 2.530 ;
        RECT 423.265 1.850 423.595 1.865 ;
        RECT 423.265 1.550 438.530 1.850 ;
        RECT 423.265 1.535 423.595 1.550 ;
        RECT 438.230 1.170 438.530 1.550 ;
        RECT 494.350 1.170 494.650 2.215 ;
        RECT 438.230 0.870 494.650 1.170 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.530 14.010 510.670 15.300 ;
        RECT 510.300 13.870 510.670 14.010 ;
        RECT 510.300 3.925 510.440 13.870 ;
        RECT 510.230 3.555 510.510 3.925 ;
        RECT 438.930 1.770 439.210 1.885 ;
        RECT 439.710 1.770 440.270 2.400 ;
        RECT 438.930 1.630 440.270 1.770 ;
        RECT 438.930 1.515 439.210 1.630 ;
        RECT 439.710 -4.800 440.270 1.630 ;
      LAYER met3 ;
        RECT 510.205 3.890 510.535 3.905 ;
        RECT 489.750 3.590 510.535 3.890 ;
        RECT 438.905 1.850 439.235 1.865 ;
        RECT 489.750 1.850 490.050 3.590 ;
        RECT 510.205 3.575 510.535 3.590 ;
        RECT 438.905 1.550 490.050 1.850 ;
        RECT 438.905 1.535 439.235 1.550 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.090 14.125 527.230 15.300 ;
        RECT 457.790 13.755 458.070 14.125 ;
        RECT 527.020 13.755 527.300 14.125 ;
        RECT 457.860 2.400 458.000 13.755 ;
        RECT 457.650 -4.800 458.210 2.400 ;
      LAYER met3 ;
        RECT 457.765 14.090 458.095 14.105 ;
        RECT 526.995 14.090 527.325 14.105 ;
        RECT 457.765 13.790 527.325 14.090 ;
        RECT 457.765 13.775 458.095 13.790 ;
        RECT 526.995 13.775 527.325 13.790 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.790 1.600 475.110 1.660 ;
        RECT 543.330 1.600 543.650 1.660 ;
        RECT 474.790 1.460 543.650 1.600 ;
        RECT 474.790 1.400 475.110 1.460 ;
        RECT 543.330 1.400 543.650 1.460 ;
      LAYER met2 ;
        RECT 543.650 14.010 543.790 15.300 ;
        RECT 543.420 13.870 543.790 14.010 ;
        RECT 475.590 1.770 476.150 2.400 ;
        RECT 474.880 1.690 476.150 1.770 ;
        RECT 543.420 1.690 543.560 13.870 ;
        RECT 474.820 1.630 476.150 1.690 ;
        RECT 474.820 1.370 475.080 1.630 ;
        RECT 475.590 -4.800 476.150 1.630 ;
        RECT 543.360 1.370 543.620 1.690 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 493.190 3.300 493.510 3.360 ;
        RECT 559.890 3.300 560.210 3.360 ;
        RECT 493.190 3.160 560.210 3.300 ;
        RECT 493.190 3.100 493.510 3.160 ;
        RECT 559.890 3.100 560.210 3.160 ;
      LAYER met2 ;
        RECT 560.210 14.010 560.350 15.300 ;
        RECT 559.980 13.870 560.350 14.010 ;
        RECT 559.980 3.390 560.120 13.870 ;
        RECT 493.220 3.070 493.480 3.390 ;
        RECT 559.920 3.070 560.180 3.390 ;
        RECT 493.280 2.400 493.420 3.070 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.770 14.010 576.910 15.300 ;
        RECT 576.540 13.870 576.910 14.010 ;
        RECT 576.540 12.085 576.680 13.870 ;
        RECT 511.150 11.715 511.430 12.085 ;
        RECT 576.470 11.715 576.750 12.085 ;
        RECT 511.220 2.400 511.360 11.715 ;
        RECT 511.010 -4.800 511.570 2.400 ;
      LAYER met3 ;
        RECT 511.125 12.050 511.455 12.065 ;
        RECT 576.445 12.050 576.775 12.065 ;
        RECT 511.125 11.750 576.775 12.050 ;
        RECT 511.125 11.735 511.455 11.750 ;
        RECT 576.445 11.735 576.775 11.750 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.330 14.010 593.470 15.300 ;
        RECT 593.100 13.870 593.470 14.010 ;
        RECT 593.100 12.765 593.240 13.870 ;
        RECT 528.630 12.395 528.910 12.765 ;
        RECT 593.030 12.395 593.310 12.765 ;
        RECT 528.700 2.400 528.840 12.395 ;
        RECT 528.490 -4.800 529.050 2.400 ;
      LAYER met3 ;
        RECT 528.605 12.730 528.935 12.745 ;
        RECT 593.005 12.730 593.335 12.745 ;
        RECT 528.605 12.430 593.335 12.730 ;
        RECT 528.605 12.415 528.935 12.430 ;
        RECT 593.005 12.415 593.335 12.430 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.890 14.010 610.030 15.300 ;
        RECT 609.660 13.870 610.030 14.010 ;
        RECT 609.660 13.445 609.800 13.870 ;
        RECT 546.570 13.075 546.850 13.445 ;
        RECT 609.590 13.075 609.870 13.445 ;
        RECT 546.640 2.400 546.780 13.075 ;
        RECT 546.430 -4.800 546.990 2.400 ;
      LAYER met3 ;
        RECT 546.545 13.410 546.875 13.425 ;
        RECT 609.565 13.410 609.895 13.425 ;
        RECT 546.545 13.110 609.895 13.410 ;
        RECT 546.545 13.095 546.875 13.110 ;
        RECT 609.565 13.095 609.895 13.110 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.450 14.010 626.590 15.300 ;
        RECT 626.220 13.870 626.590 14.010 ;
        RECT 626.220 8.685 626.360 13.870 ;
        RECT 564.050 8.315 564.330 8.685 ;
        RECT 626.150 8.315 626.430 8.685 ;
        RECT 564.120 2.400 564.260 8.315 ;
        RECT 563.910 -4.800 564.470 2.400 ;
      LAYER met3 ;
        RECT 564.025 8.650 564.355 8.665 ;
        RECT 626.125 8.650 626.455 8.665 ;
        RECT 564.025 8.350 626.455 8.650 ;
        RECT 564.025 8.335 564.355 8.350 ;
        RECT 626.125 8.335 626.455 8.350 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.430 6.020 582.750 6.080 ;
        RECT 642.690 6.020 643.010 6.080 ;
        RECT 582.430 5.880 643.010 6.020 ;
        RECT 582.430 5.820 582.750 5.880 ;
        RECT 642.690 5.820 643.010 5.880 ;
      LAYER met2 ;
        RECT 643.010 14.010 643.150 15.300 ;
        RECT 642.780 13.870 643.150 14.010 ;
        RECT 642.780 6.110 642.920 13.870 ;
        RECT 582.460 5.790 582.720 6.110 ;
        RECT 642.720 5.790 642.980 6.110 ;
        RECT 582.520 3.130 582.660 5.790 ;
        RECT 582.060 2.990 582.660 3.130 ;
        RECT 582.060 2.400 582.200 2.990 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.850 14.010 184.990 15.300 ;
        RECT 184.620 13.870 184.990 14.010 ;
        RECT 184.620 3.925 184.760 13.870 ;
        RECT 91.170 3.555 91.450 3.925 ;
        RECT 184.550 3.555 184.830 3.925 ;
        RECT 91.240 2.400 91.380 3.555 ;
        RECT 91.030 -4.800 91.590 2.400 ;
      LAYER met3 ;
        RECT 91.145 3.890 91.475 3.905 ;
        RECT 184.525 3.890 184.855 3.905 ;
        RECT 91.145 3.590 184.855 3.890 ;
        RECT 91.145 3.575 91.475 3.590 ;
        RECT 184.525 3.575 184.855 3.590 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 659.250 7.040 659.570 7.100 ;
        RECT 657.960 6.900 659.570 7.040 ;
        RECT 599.450 6.700 599.770 6.760 ;
        RECT 657.960 6.700 658.100 6.900 ;
        RECT 659.250 6.840 659.570 6.900 ;
        RECT 599.450 6.560 658.100 6.700 ;
        RECT 599.450 6.500 599.770 6.560 ;
      LAYER met2 ;
        RECT 659.570 14.010 659.710 15.300 ;
        RECT 659.340 13.870 659.710 14.010 ;
        RECT 659.340 7.130 659.480 13.870 ;
        RECT 659.280 6.810 659.540 7.130 ;
        RECT 599.480 6.470 599.740 6.790 ;
        RECT 599.540 2.400 599.680 6.470 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.130 14.010 676.270 15.300 ;
        RECT 675.900 13.870 676.270 14.010 ;
        RECT 675.900 3.925 676.040 13.870 ;
        RECT 617.410 3.555 617.690 3.925 ;
        RECT 675.830 3.555 676.110 3.925 ;
        RECT 617.480 2.400 617.620 3.555 ;
        RECT 617.270 -4.800 617.830 2.400 ;
      LAYER met3 ;
        RECT 617.385 3.890 617.715 3.905 ;
        RECT 675.805 3.890 676.135 3.905 ;
        RECT 617.385 3.590 676.135 3.890 ;
        RECT 617.385 3.575 617.715 3.590 ;
        RECT 675.805 3.575 676.135 3.590 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.930 14.125 207.070 15.300 ;
        RECT 115.090 13.755 115.370 14.125 ;
        RECT 206.860 13.755 207.140 14.125 ;
        RECT 115.160 2.400 115.300 13.755 ;
        RECT 114.950 -4.800 115.510 2.400 ;
      LAYER met3 ;
        RECT 115.065 14.090 115.395 14.105 ;
        RECT 206.835 14.090 207.165 14.105 ;
        RECT 115.065 13.790 207.165 14.090 ;
        RECT 115.065 13.775 115.395 13.790 ;
        RECT 206.835 13.775 207.165 13.790 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 184.990 5.340 185.310 5.400 ;
        RECT 228.690 5.340 229.010 5.400 ;
        RECT 184.990 5.200 229.010 5.340 ;
        RECT 184.990 5.140 185.310 5.200 ;
        RECT 228.690 5.140 229.010 5.200 ;
      LAYER met2 ;
        RECT 229.010 14.010 229.150 15.300 ;
        RECT 228.780 13.870 229.150 14.010 ;
        RECT 228.780 5.430 228.920 13.870 ;
        RECT 185.020 5.110 185.280 5.430 ;
        RECT 228.720 5.110 228.980 5.430 ;
        RECT 185.080 2.565 185.220 5.110 ;
        RECT 138.410 1.770 138.970 2.400 ;
        RECT 140.850 2.195 141.130 2.565 ;
        RECT 185.010 2.195 185.290 2.565 ;
        RECT 140.920 1.770 141.060 2.195 ;
        RECT 138.410 1.630 141.060 1.770 ;
        RECT 138.410 -4.800 138.970 1.630 ;
      LAYER met3 ;
        RECT 140.825 2.530 141.155 2.545 ;
        RECT 184.985 2.530 185.315 2.545 ;
        RECT 140.825 2.230 185.315 2.530 ;
        RECT 140.825 2.215 141.155 2.230 ;
        RECT 184.985 2.215 185.315 2.230 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 166.130 5.000 166.450 5.060 ;
        RECT 245.250 5.000 245.570 5.060 ;
        RECT 166.130 4.860 245.570 5.000 ;
        RECT 166.130 4.800 166.450 4.860 ;
        RECT 245.250 4.800 245.570 4.860 ;
      LAYER met2 ;
        RECT 245.570 14.010 245.710 15.300 ;
        RECT 245.340 13.870 245.710 14.010 ;
        RECT 245.340 5.090 245.480 13.870 ;
        RECT 166.160 4.770 166.420 5.090 ;
        RECT 245.280 4.770 245.540 5.090 ;
        RECT 166.220 3.245 166.360 4.770 ;
        RECT 156.490 2.875 156.770 3.245 ;
        RECT 166.150 2.875 166.430 3.245 ;
        RECT 156.560 2.400 156.700 2.875 ;
        RECT 156.350 -4.800 156.910 2.400 ;
      LAYER met3 ;
        RECT 156.465 3.210 156.795 3.225 ;
        RECT 166.125 3.210 166.455 3.225 ;
        RECT 156.465 2.910 166.455 3.210 ;
        RECT 156.465 2.895 156.795 2.910 ;
        RECT 166.125 2.895 166.455 2.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.130 14.805 262.270 15.300 ;
        RECT 262.060 14.435 262.340 14.805 ;
        RECT 173.970 12.395 174.250 12.765 ;
        RECT 174.040 2.400 174.180 12.395 ;
        RECT 173.830 -4.800 174.390 2.400 ;
      LAYER met3 ;
        RECT 174.150 16.130 174.530 16.140 ;
        RECT 174.150 15.830 227.850 16.130 ;
        RECT 174.150 15.820 174.530 15.830 ;
        RECT 227.550 14.770 227.850 15.830 ;
        RECT 262.035 14.770 262.365 14.785 ;
        RECT 227.550 14.470 262.365 14.770 ;
        RECT 262.035 14.455 262.365 14.470 ;
        RECT 173.945 12.740 174.275 12.745 ;
        RECT 173.945 12.730 174.530 12.740 ;
        RECT 173.720 12.430 174.530 12.730 ;
        RECT 173.945 12.420 174.530 12.430 ;
        RECT 173.945 12.415 174.275 12.420 ;
      LAYER met4 ;
        RECT 174.175 15.815 174.505 16.145 ;
        RECT 174.190 12.745 174.490 15.815 ;
        RECT 174.175 12.415 174.505 12.745 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.810 1.260 193.130 1.320 ;
        RECT 278.370 1.260 278.690 1.320 ;
        RECT 192.810 1.120 278.690 1.260 ;
        RECT 192.810 1.060 193.130 1.120 ;
        RECT 278.370 1.060 278.690 1.120 ;
      LAYER met2 ;
        RECT 278.690 14.010 278.830 15.300 ;
        RECT 278.460 13.870 278.830 14.010 ;
        RECT 191.770 1.090 192.330 2.400 ;
        RECT 278.460 1.350 278.600 13.870 ;
        RECT 192.840 1.090 193.100 1.350 ;
        RECT 191.770 1.030 193.100 1.090 ;
        RECT 278.400 1.030 278.660 1.350 ;
        RECT 191.770 0.950 193.040 1.030 ;
        RECT 191.770 -4.800 192.330 0.950 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 209.370 14.180 209.690 14.240 ;
        RECT 248.010 14.180 248.330 14.240 ;
        RECT 209.370 14.040 248.330 14.180 ;
        RECT 209.370 13.980 209.690 14.040 ;
        RECT 248.010 13.980 248.330 14.040 ;
        RECT 248.010 6.360 248.330 6.420 ;
        RECT 294.930 6.360 295.250 6.420 ;
        RECT 248.010 6.220 295.250 6.360 ;
        RECT 248.010 6.160 248.330 6.220 ;
        RECT 294.930 6.160 295.250 6.220 ;
      LAYER met2 ;
        RECT 209.400 13.950 209.660 14.270 ;
        RECT 248.040 13.950 248.300 14.270 ;
        RECT 295.250 14.010 295.390 15.300 ;
        RECT 209.460 2.400 209.600 13.950 ;
        RECT 248.100 6.450 248.240 13.950 ;
        RECT 295.020 13.870 295.390 14.010 ;
        RECT 295.020 6.450 295.160 13.870 ;
        RECT 248.040 6.130 248.300 6.450 ;
        RECT 294.960 6.130 295.220 6.450 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 227.310 2.960 227.630 3.020 ;
        RECT 311.490 2.960 311.810 3.020 ;
        RECT 227.310 2.820 311.810 2.960 ;
        RECT 227.310 2.760 227.630 2.820 ;
        RECT 311.490 2.760 311.810 2.820 ;
      LAYER met2 ;
        RECT 311.810 14.010 311.950 15.300 ;
        RECT 311.580 13.870 311.950 14.010 ;
        RECT 311.580 3.050 311.720 13.870 ;
        RECT 227.340 2.730 227.600 3.050 ;
        RECT 311.520 2.730 311.780 3.050 ;
        RECT 227.400 2.400 227.540 2.730 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 49.750 4.320 50.070 4.380 ;
        RECT 145.890 4.320 146.210 4.380 ;
        RECT 49.750 4.180 146.210 4.320 ;
        RECT 49.750 4.120 50.070 4.180 ;
        RECT 145.890 4.120 146.210 4.180 ;
      LAYER met2 ;
        RECT 146.210 14.010 146.350 15.300 ;
        RECT 145.980 13.870 146.350 14.010 ;
        RECT 145.980 4.410 146.120 13.870 ;
        RECT 49.780 4.090 50.040 4.410 ;
        RECT 145.920 4.090 146.180 4.410 ;
        RECT 49.840 2.400 49.980 4.090 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 250.770 3.640 251.090 3.700 ;
        RECT 333.570 3.640 333.890 3.700 ;
        RECT 250.770 3.500 333.890 3.640 ;
        RECT 250.770 3.440 251.090 3.500 ;
        RECT 333.570 3.440 333.890 3.500 ;
      LAYER met2 ;
        RECT 333.890 14.010 334.030 15.300 ;
        RECT 333.660 13.870 334.030 14.010 ;
        RECT 333.660 3.730 333.800 13.870 ;
        RECT 250.800 3.410 251.060 3.730 ;
        RECT 333.600 3.410 333.860 3.730 ;
        RECT 250.860 2.400 251.000 3.410 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 267.790 0.580 268.110 0.640 ;
        RECT 350.130 0.580 350.450 0.640 ;
        RECT 267.790 0.440 350.450 0.580 ;
        RECT 267.790 0.380 268.110 0.440 ;
        RECT 350.130 0.380 350.450 0.440 ;
      LAYER met2 ;
        RECT 350.450 14.010 350.590 15.300 ;
        RECT 350.220 13.870 350.590 14.010 ;
        RECT 267.820 0.410 268.080 0.670 ;
        RECT 268.590 0.410 269.150 2.400 ;
        RECT 350.220 0.670 350.360 13.870 ;
        RECT 267.820 0.350 269.150 0.410 ;
        RECT 350.160 0.350 350.420 0.670 ;
        RECT 267.880 0.270 269.150 0.350 ;
        RECT 268.590 -4.800 269.150 0.270 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 285.270 1.600 285.590 1.660 ;
        RECT 366.690 1.600 367.010 1.660 ;
        RECT 285.270 1.460 367.010 1.600 ;
        RECT 285.270 1.400 285.590 1.460 ;
        RECT 366.690 1.400 367.010 1.460 ;
      LAYER met2 ;
        RECT 367.010 14.010 367.150 15.300 ;
        RECT 366.780 13.870 367.150 14.010 ;
        RECT 286.070 1.770 286.630 2.400 ;
        RECT 285.360 1.690 286.630 1.770 ;
        RECT 366.780 1.690 366.920 13.870 ;
        RECT 285.300 1.630 286.630 1.690 ;
        RECT 285.300 1.370 285.560 1.630 ;
        RECT 286.070 -4.800 286.630 1.630 ;
        RECT 366.720 1.370 366.980 1.690 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.130 14.180 304.450 14.240 ;
        RECT 344.610 14.180 344.930 14.240 ;
        RECT 304.130 14.040 344.930 14.180 ;
        RECT 304.130 13.980 304.450 14.040 ;
        RECT 344.610 13.980 344.930 14.040 ;
        RECT 344.610 6.700 344.930 6.760 ;
        RECT 383.250 6.700 383.570 6.760 ;
        RECT 344.610 6.560 383.570 6.700 ;
        RECT 344.610 6.500 344.930 6.560 ;
        RECT 383.250 6.500 383.570 6.560 ;
      LAYER met2 ;
        RECT 304.160 13.950 304.420 14.270 ;
        RECT 344.640 13.950 344.900 14.270 ;
        RECT 383.570 14.010 383.710 15.300 ;
        RECT 304.220 2.400 304.360 13.950 ;
        RECT 344.700 6.790 344.840 13.950 ;
        RECT 383.340 13.870 383.710 14.010 ;
        RECT 383.340 6.790 383.480 13.870 ;
        RECT 344.640 6.470 344.900 6.790 ;
        RECT 383.280 6.470 383.540 6.790 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 321.610 2.960 321.930 3.020 ;
        RECT 399.810 2.960 400.130 3.020 ;
        RECT 321.610 2.820 400.130 2.960 ;
        RECT 321.610 2.760 321.930 2.820 ;
        RECT 399.810 2.760 400.130 2.820 ;
      LAYER met2 ;
        RECT 400.130 14.010 400.270 15.300 ;
        RECT 399.900 13.870 400.270 14.010 ;
        RECT 399.900 3.050 400.040 13.870 ;
        RECT 321.640 2.730 321.900 3.050 ;
        RECT 399.840 2.730 400.100 3.050 ;
        RECT 321.700 2.400 321.840 2.730 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 416.370 6.700 416.690 6.760 ;
        RECT 385.640 6.560 416.690 6.700 ;
        RECT 339.550 6.020 339.870 6.080 ;
        RECT 385.640 6.020 385.780 6.560 ;
        RECT 416.370 6.500 416.690 6.560 ;
        RECT 339.550 5.880 385.780 6.020 ;
        RECT 339.550 5.820 339.870 5.880 ;
      LAYER met2 ;
        RECT 416.690 14.010 416.830 15.300 ;
        RECT 416.460 13.870 416.830 14.010 ;
        RECT 416.460 6.790 416.600 13.870 ;
        RECT 416.400 6.470 416.660 6.790 ;
        RECT 339.580 5.790 339.840 6.110 ;
        RECT 339.640 2.400 339.780 5.790 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.410 0.580 358.730 0.640 ;
        RECT 432.930 0.580 433.250 0.640 ;
        RECT 358.410 0.440 433.250 0.580 ;
        RECT 358.410 0.380 358.730 0.440 ;
        RECT 432.930 0.380 433.250 0.440 ;
      LAYER met2 ;
        RECT 433.250 14.010 433.390 15.300 ;
        RECT 433.020 13.870 433.390 14.010 ;
        RECT 357.370 0.410 357.930 2.400 ;
        RECT 433.020 0.670 433.160 13.870 ;
        RECT 358.440 0.410 358.700 0.670 ;
        RECT 357.370 0.350 358.700 0.410 ;
        RECT 432.960 0.350 433.220 0.670 ;
        RECT 357.370 0.270 358.640 0.350 ;
        RECT 357.370 -4.800 357.930 0.270 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 376.810 1.260 377.130 1.320 ;
        RECT 449.490 1.260 449.810 1.320 ;
        RECT 376.810 1.120 449.810 1.260 ;
        RECT 376.810 1.060 377.130 1.120 ;
        RECT 449.490 1.060 449.810 1.120 ;
      LAYER met2 ;
        RECT 449.810 14.010 449.950 15.300 ;
        RECT 449.580 13.870 449.950 14.010 ;
        RECT 374.850 1.090 375.410 2.400 ;
        RECT 449.580 1.350 449.720 13.870 ;
        RECT 376.840 1.090 377.100 1.350 ;
        RECT 374.850 1.030 377.100 1.090 ;
        RECT 449.520 1.030 449.780 1.350 ;
        RECT 374.850 0.950 377.040 1.030 ;
        RECT 374.850 -4.800 375.410 0.950 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 391.990 1.940 392.310 2.000 ;
        RECT 466.050 1.940 466.370 2.000 ;
        RECT 391.990 1.800 466.370 1.940 ;
        RECT 391.990 1.740 392.310 1.800 ;
        RECT 466.050 1.740 466.370 1.800 ;
      LAYER met2 ;
        RECT 466.370 14.010 466.510 15.300 ;
        RECT 466.140 13.870 466.510 14.010 ;
        RECT 392.020 1.770 392.280 2.030 ;
        RECT 392.790 1.770 393.350 2.400 ;
        RECT 466.140 2.030 466.280 13.870 ;
        RECT 392.020 1.710 393.350 1.770 ;
        RECT 466.080 1.710 466.340 2.030 ;
        RECT 392.080 1.630 393.350 1.710 ;
        RECT 392.790 -4.800 393.350 1.630 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 410.390 14.180 410.710 14.240 ;
        RECT 482.840 14.180 483.160 14.240 ;
        RECT 410.390 14.040 483.160 14.180 ;
        RECT 410.390 13.980 410.710 14.040 ;
        RECT 482.840 13.980 483.160 14.040 ;
      LAYER met2 ;
        RECT 482.930 14.270 483.070 15.300 ;
        RECT 410.420 13.950 410.680 14.270 ;
        RECT 482.870 13.950 483.130 14.270 ;
        RECT 410.480 2.400 410.620 13.950 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 72.750 0.920 73.070 0.980 ;
        RECT 167.050 0.920 167.370 0.980 ;
        RECT 72.750 0.780 167.370 0.920 ;
        RECT 72.750 0.720 73.070 0.780 ;
        RECT 167.050 0.720 167.370 0.780 ;
      LAYER met2 ;
        RECT 168.290 14.010 168.430 15.300 ;
        RECT 167.140 13.870 168.430 14.010 ;
        RECT 73.550 1.090 74.110 2.400 ;
        RECT 72.840 1.010 74.110 1.090 ;
        RECT 167.140 1.010 167.280 13.870 ;
        RECT 72.780 0.950 74.110 1.010 ;
        RECT 72.780 0.690 73.040 0.950 ;
        RECT 73.550 -4.800 74.110 0.950 ;
        RECT 167.080 0.690 167.340 1.010 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 499.630 2.760 499.950 3.020 ;
        RECT 430.630 2.280 430.950 2.340 ;
        RECT 499.720 2.280 499.860 2.760 ;
        RECT 430.630 2.140 499.860 2.280 ;
        RECT 430.630 2.080 430.950 2.140 ;
      LAYER met2 ;
        RECT 499.490 14.010 499.630 15.300 ;
        RECT 499.490 13.870 499.860 14.010 ;
        RECT 499.720 3.050 499.860 13.870 ;
        RECT 499.660 2.730 499.920 3.050 ;
        RECT 428.210 1.770 428.770 2.400 ;
        RECT 430.660 2.050 430.920 2.370 ;
        RECT 430.720 1.770 430.860 2.050 ;
        RECT 428.210 1.630 430.860 1.770 ;
        RECT 428.210 -4.800 428.770 1.630 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 447.650 0.920 447.970 0.980 ;
        RECT 515.730 0.920 516.050 0.980 ;
        RECT 447.650 0.780 516.050 0.920 ;
        RECT 447.650 0.720 447.970 0.780 ;
        RECT 515.730 0.720 516.050 0.780 ;
      LAYER met2 ;
        RECT 516.050 14.010 516.190 15.300 ;
        RECT 515.820 13.870 516.190 14.010 ;
        RECT 445.690 1.090 446.250 2.400 ;
        RECT 445.690 1.010 447.880 1.090 ;
        RECT 515.820 1.010 515.960 13.870 ;
        RECT 445.690 0.950 447.940 1.010 ;
        RECT 445.690 -4.800 446.250 0.950 ;
        RECT 447.680 0.690 447.940 0.950 ;
        RECT 515.760 0.690 516.020 1.010 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.830 1.260 463.150 1.320 ;
        RECT 532.290 1.260 532.610 1.320 ;
        RECT 462.830 1.120 532.610 1.260 ;
        RECT 462.830 1.060 463.150 1.120 ;
        RECT 532.290 1.060 532.610 1.120 ;
      LAYER met2 ;
        RECT 532.610 14.010 532.750 15.300 ;
        RECT 532.380 13.870 532.750 14.010 ;
        RECT 462.860 1.090 463.120 1.350 ;
        RECT 463.630 1.090 464.190 2.400 ;
        RECT 532.380 1.350 532.520 13.870 ;
        RECT 462.860 1.030 464.190 1.090 ;
        RECT 532.320 1.030 532.580 1.350 ;
        RECT 462.920 0.950 464.190 1.030 ;
        RECT 463.630 -4.800 464.190 0.950 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 480.310 1.940 480.630 2.000 ;
        RECT 548.850 1.940 549.170 2.000 ;
        RECT 480.310 1.800 549.170 1.940 ;
        RECT 480.310 1.740 480.630 1.800 ;
        RECT 548.850 1.740 549.170 1.800 ;
      LAYER met2 ;
        RECT 549.170 14.010 549.310 15.300 ;
        RECT 548.940 13.870 549.310 14.010 ;
        RECT 480.340 1.770 480.600 2.030 ;
        RECT 481.110 1.770 481.670 2.400 ;
        RECT 548.940 2.030 549.080 13.870 ;
        RECT 480.340 1.710 481.670 1.770 ;
        RECT 548.880 1.710 549.140 2.030 ;
        RECT 480.400 1.630 481.670 1.710 ;
        RECT 481.110 -4.800 481.670 1.630 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.730 14.010 565.870 15.300 ;
        RECT 565.500 13.870 565.870 14.010 ;
        RECT 565.500 11.405 565.640 13.870 ;
        RECT 498.730 11.035 499.010 11.405 ;
        RECT 565.430 11.035 565.710 11.405 ;
        RECT 498.800 3.130 498.940 11.035 ;
        RECT 498.800 2.990 499.400 3.130 ;
        RECT 499.260 2.400 499.400 2.990 ;
        RECT 499.050 -4.800 499.610 2.400 ;
      LAYER met3 ;
        RECT 498.705 11.370 499.035 11.385 ;
        RECT 565.405 11.370 565.735 11.385 ;
        RECT 498.705 11.070 565.735 11.370 ;
        RECT 498.705 11.055 499.035 11.070 ;
        RECT 565.405 11.055 565.735 11.070 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 0.580 517.890 0.640 ;
        RECT 581.050 0.580 581.370 0.640 ;
        RECT 517.570 0.440 581.370 0.580 ;
        RECT 517.570 0.380 517.890 0.440 ;
        RECT 581.050 0.380 581.370 0.440 ;
      LAYER met2 ;
        RECT 582.290 14.010 582.430 15.300 ;
        RECT 581.140 13.870 582.430 14.010 ;
        RECT 516.530 0.410 517.090 2.400 ;
        RECT 581.140 0.670 581.280 13.870 ;
        RECT 517.600 0.410 517.860 0.670 ;
        RECT 516.530 0.350 517.860 0.410 ;
        RECT 581.080 0.350 581.340 0.670 ;
        RECT 516.530 0.270 517.800 0.350 ;
        RECT 516.530 -4.800 517.090 0.270 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.970 6.360 536.290 6.420 ;
        RECT 598.530 6.360 598.850 6.420 ;
        RECT 535.970 6.220 598.850 6.360 ;
        RECT 535.970 6.160 536.290 6.220 ;
        RECT 598.530 6.160 598.850 6.220 ;
      LAYER met2 ;
        RECT 598.850 14.010 598.990 15.300 ;
        RECT 598.620 13.870 598.990 14.010 ;
        RECT 598.620 6.450 598.760 13.870 ;
        RECT 536.000 6.130 536.260 6.450 ;
        RECT 598.560 6.130 598.820 6.450 ;
        RECT 536.060 3.130 536.200 6.130 ;
        RECT 534.680 2.990 536.200 3.130 ;
        RECT 534.680 2.400 534.820 2.990 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.830 5.680 555.150 5.740 ;
        RECT 615.090 5.680 615.410 5.740 ;
        RECT 554.830 5.540 615.410 5.680 ;
        RECT 554.830 5.480 555.150 5.540 ;
        RECT 615.090 5.480 615.410 5.540 ;
      LAYER met2 ;
        RECT 615.410 14.010 615.550 15.300 ;
        RECT 615.180 13.870 615.550 14.010 ;
        RECT 615.180 5.770 615.320 13.870 ;
        RECT 554.860 5.450 555.120 5.770 ;
        RECT 615.120 5.450 615.380 5.770 ;
        RECT 552.410 1.770 552.970 2.400 ;
        RECT 554.920 1.770 555.060 5.450 ;
        RECT 552.410 1.630 555.060 1.770 ;
        RECT 552.410 -4.800 552.970 1.630 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.850 0.920 572.170 0.980 ;
        RECT 631.650 0.920 631.970 0.980 ;
        RECT 571.850 0.780 631.970 0.920 ;
        RECT 571.850 0.720 572.170 0.780 ;
        RECT 631.650 0.720 631.970 0.780 ;
      LAYER met2 ;
        RECT 631.970 14.010 632.110 15.300 ;
        RECT 631.740 13.870 632.110 14.010 ;
        RECT 569.890 1.090 570.450 2.400 ;
        RECT 569.890 1.010 572.080 1.090 ;
        RECT 631.740 1.010 631.880 13.870 ;
        RECT 569.890 0.950 572.140 1.010 ;
        RECT 569.890 -4.800 570.450 0.950 ;
        RECT 571.880 0.690 572.140 0.950 ;
        RECT 631.680 0.690 631.940 1.010 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.530 14.125 648.670 15.300 ;
        RECT 588.430 13.755 588.710 14.125 ;
        RECT 648.460 13.755 648.740 14.125 ;
        RECT 588.500 7.210 588.640 13.755 ;
        RECT 588.040 7.070 588.640 7.210 ;
        RECT 588.040 2.400 588.180 7.070 ;
        RECT 587.830 -4.800 588.390 2.400 ;
      LAYER met3 ;
        RECT 588.405 14.090 588.735 14.105 ;
        RECT 648.435 14.090 648.765 14.105 ;
        RECT 588.405 13.790 648.765 14.090 ;
        RECT 588.405 13.775 588.735 13.790 ;
        RECT 648.435 13.775 648.765 13.790 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 155.090 6.700 155.410 6.760 ;
        RECT 190.050 6.700 190.370 6.760 ;
        RECT 155.090 6.560 190.370 6.700 ;
        RECT 155.090 6.500 155.410 6.560 ;
        RECT 190.050 6.500 190.370 6.560 ;
      LAYER met2 ;
        RECT 190.370 14.010 190.510 15.300 ;
        RECT 190.140 13.870 190.510 14.010 ;
        RECT 190.140 6.790 190.280 13.870 ;
        RECT 155.120 6.470 155.380 6.790 ;
        RECT 190.080 6.470 190.340 6.790 ;
        RECT 155.180 4.605 155.320 6.470 ;
        RECT 97.150 4.235 97.430 4.605 ;
        RECT 155.110 4.235 155.390 4.605 ;
        RECT 97.220 2.400 97.360 4.235 ;
        RECT 97.010 -4.800 97.570 2.400 ;
      LAYER met3 ;
        RECT 97.125 4.570 97.455 4.585 ;
        RECT 155.085 4.570 155.415 4.585 ;
        RECT 97.125 4.270 155.415 4.570 ;
        RECT 97.125 4.255 97.455 4.270 ;
        RECT 155.085 4.255 155.415 4.270 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.810 6.360 607.130 6.420 ;
        RECT 664.770 6.360 665.090 6.420 ;
        RECT 606.810 6.220 665.090 6.360 ;
        RECT 606.810 6.160 607.130 6.220 ;
        RECT 664.770 6.160 665.090 6.220 ;
      LAYER met2 ;
        RECT 665.090 14.010 665.230 15.300 ;
        RECT 664.860 13.870 665.230 14.010 ;
        RECT 664.860 6.450 665.000 13.870 ;
        RECT 606.840 6.130 607.100 6.450 ;
        RECT 664.800 6.130 665.060 6.450 ;
        RECT 606.900 3.130 607.040 6.130 ;
        RECT 605.520 2.990 607.040 3.130 ;
        RECT 605.520 2.400 605.660 2.990 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 681.330 6.020 681.650 6.080 ;
        RECT 662.330 5.880 681.650 6.020 ;
        RECT 625.670 5.680 625.990 5.740 ;
        RECT 662.330 5.680 662.470 5.880 ;
        RECT 681.330 5.820 681.650 5.880 ;
        RECT 625.670 5.540 662.470 5.680 ;
        RECT 625.670 5.480 625.990 5.540 ;
      LAYER met2 ;
        RECT 681.650 14.010 681.790 15.300 ;
        RECT 681.420 13.870 681.790 14.010 ;
        RECT 681.420 6.110 681.560 13.870 ;
        RECT 681.360 5.790 681.620 6.110 ;
        RECT 625.700 5.450 625.960 5.770 ;
        RECT 623.250 1.770 623.810 2.400 ;
        RECT 625.760 1.770 625.900 5.450 ;
        RECT 623.250 1.630 625.900 1.770 ;
        RECT 623.250 -4.800 623.810 1.630 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 151.410 5.680 151.730 5.740 ;
        RECT 212.130 5.680 212.450 5.740 ;
        RECT 151.410 5.540 212.450 5.680 ;
        RECT 151.410 5.480 151.730 5.540 ;
        RECT 212.130 5.480 212.450 5.540 ;
      LAYER met2 ;
        RECT 212.450 14.010 212.590 15.300 ;
        RECT 212.220 13.870 212.590 14.010 ;
        RECT 212.220 5.770 212.360 13.870 ;
        RECT 151.440 5.450 151.700 5.770 ;
        RECT 212.160 5.450 212.420 5.770 ;
        RECT 120.930 1.770 121.490 2.400 ;
        RECT 151.500 1.885 151.640 5.450 ;
        RECT 123.830 1.770 124.110 1.885 ;
        RECT 120.930 1.630 124.110 1.770 ;
        RECT 120.930 -4.800 121.490 1.630 ;
        RECT 123.830 1.515 124.110 1.630 ;
        RECT 151.430 1.515 151.710 1.885 ;
      LAYER met3 ;
        RECT 123.805 1.850 124.135 1.865 ;
        RECT 151.405 1.850 151.735 1.865 ;
        RECT 123.805 1.550 151.735 1.850 ;
        RECT 123.805 1.535 124.135 1.550 ;
        RECT 151.405 1.535 151.735 1.550 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 143.590 1.940 143.910 2.000 ;
        RECT 234.210 1.940 234.530 2.000 ;
        RECT 143.590 1.800 234.530 1.940 ;
        RECT 143.590 1.740 143.910 1.800 ;
        RECT 234.210 1.740 234.530 1.800 ;
      LAYER met2 ;
        RECT 234.530 14.010 234.670 15.300 ;
        RECT 234.300 13.870 234.670 14.010 ;
        RECT 143.620 1.770 143.880 2.030 ;
        RECT 144.390 1.770 144.950 2.400 ;
        RECT 234.300 2.030 234.440 13.870 ;
        RECT 143.620 1.710 144.950 1.770 ;
        RECT 234.240 1.710 234.500 2.030 ;
        RECT 143.680 1.630 144.950 1.710 ;
        RECT 144.390 -4.800 144.950 1.630 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.070 2.280 161.390 2.340 ;
        RECT 249.850 2.280 250.170 2.340 ;
        RECT 161.070 2.140 250.170 2.280 ;
        RECT 161.070 2.080 161.390 2.140 ;
        RECT 249.850 2.080 250.170 2.140 ;
      LAYER met2 ;
        RECT 251.090 14.010 251.230 15.300 ;
        RECT 249.940 13.870 251.230 14.010 ;
        RECT 161.100 2.050 161.360 2.370 ;
        RECT 161.160 1.770 161.300 2.050 ;
        RECT 161.870 1.770 162.430 2.400 ;
        RECT 249.940 2.370 250.080 13.870 ;
        RECT 249.880 2.050 250.140 2.370 ;
        RECT 161.160 1.630 162.430 1.770 ;
        RECT 161.870 -4.800 162.430 1.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 179.930 14.520 180.250 14.580 ;
        RECT 202.010 14.520 202.330 14.580 ;
        RECT 179.930 14.380 202.330 14.520 ;
        RECT 179.930 14.320 180.250 14.380 ;
        RECT 202.010 14.320 202.330 14.380 ;
        RECT 202.010 6.020 202.330 6.080 ;
        RECT 267.330 6.020 267.650 6.080 ;
        RECT 202.010 5.880 267.650 6.020 ;
        RECT 202.010 5.820 202.330 5.880 ;
        RECT 267.330 5.820 267.650 5.880 ;
      LAYER met2 ;
        RECT 179.960 14.290 180.220 14.610 ;
        RECT 202.040 14.290 202.300 14.610 ;
        RECT 180.020 2.400 180.160 14.290 ;
        RECT 202.100 6.110 202.240 14.290 ;
        RECT 267.650 14.010 267.790 15.300 ;
        RECT 267.420 13.870 267.790 14.010 ;
        RECT 267.420 6.110 267.560 13.870 ;
        RECT 202.040 5.790 202.300 6.110 ;
        RECT 267.360 5.790 267.620 6.110 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 196.950 1.600 197.270 1.660 ;
        RECT 283.890 1.600 284.210 1.660 ;
        RECT 196.950 1.460 284.210 1.600 ;
        RECT 196.950 1.400 197.270 1.460 ;
        RECT 283.890 1.400 284.210 1.460 ;
      LAYER met2 ;
        RECT 284.210 14.010 284.350 15.300 ;
        RECT 283.980 13.870 284.350 14.010 ;
        RECT 197.750 1.770 198.310 2.400 ;
        RECT 197.040 1.690 198.310 1.770 ;
        RECT 283.980 1.690 284.120 13.870 ;
        RECT 196.980 1.630 198.310 1.690 ;
        RECT 196.980 1.370 197.240 1.630 ;
        RECT 197.750 -4.800 198.310 1.630 ;
        RECT 283.920 1.370 284.180 1.690 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.430 2.620 214.750 2.680 ;
        RECT 300.450 2.620 300.770 2.680 ;
        RECT 214.430 2.480 300.770 2.620 ;
        RECT 214.430 2.420 214.750 2.480 ;
        RECT 300.450 2.420 300.770 2.480 ;
      LAYER met2 ;
        RECT 300.770 14.010 300.910 15.300 ;
        RECT 300.540 13.870 300.910 14.010 ;
        RECT 300.540 2.710 300.680 13.870 ;
        RECT 214.460 2.390 214.720 2.710 ;
        RECT 214.520 1.770 214.660 2.390 ;
        RECT 215.230 1.770 215.790 2.400 ;
        RECT 300.480 2.390 300.740 2.710 ;
        RECT 214.520 1.630 215.790 1.770 ;
        RECT 215.230 -4.800 215.790 1.630 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 233.290 3.300 233.610 3.360 ;
        RECT 317.010 3.300 317.330 3.360 ;
        RECT 233.290 3.160 317.330 3.300 ;
        RECT 233.290 3.100 233.610 3.160 ;
        RECT 317.010 3.100 317.330 3.160 ;
      LAYER met2 ;
        RECT 317.330 14.010 317.470 15.300 ;
        RECT 317.100 13.870 317.470 14.010 ;
        RECT 317.100 3.390 317.240 13.870 ;
        RECT 233.320 3.070 233.580 3.390 ;
        RECT 317.040 3.070 317.300 3.390 ;
        RECT 233.380 2.400 233.520 3.070 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 141.290 6.700 141.610 6.760 ;
        RECT 151.410 6.700 151.730 6.760 ;
        RECT 141.290 6.560 151.730 6.700 ;
        RECT 141.290 6.500 141.610 6.560 ;
        RECT 151.410 6.500 151.730 6.560 ;
      LAYER met2 ;
        RECT 151.730 14.010 151.870 15.300 ;
        RECT 151.500 13.870 151.870 14.010 ;
        RECT 151.500 6.790 151.640 13.870 ;
        RECT 141.320 6.470 141.580 6.790 ;
        RECT 151.440 6.470 151.700 6.790 ;
        RECT 141.380 3.245 141.520 6.470 ;
        RECT 55.750 2.875 56.030 3.245 ;
        RECT 141.310 2.875 141.590 3.245 ;
        RECT 55.820 2.400 55.960 2.875 ;
        RECT 55.610 -4.800 56.170 2.400 ;
      LAYER met3 ;
        RECT 55.725 3.210 56.055 3.225 ;
        RECT 141.285 3.210 141.615 3.225 ;
        RECT 55.725 2.910 141.615 3.210 ;
        RECT 55.725 2.895 56.055 2.910 ;
        RECT 141.285 2.895 141.615 2.910 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 81.030 1.260 81.350 1.320 ;
        RECT 173.030 1.260 173.350 1.320 ;
        RECT 81.030 1.120 173.350 1.260 ;
        RECT 81.030 1.060 81.350 1.120 ;
        RECT 173.030 1.060 173.350 1.120 ;
      LAYER met2 ;
        RECT 173.810 14.010 173.950 15.300 ;
        RECT 173.120 13.870 173.950 14.010 ;
        RECT 79.530 1.090 80.090 2.400 ;
        RECT 173.120 1.350 173.260 13.870 ;
        RECT 81.060 1.090 81.320 1.350 ;
        RECT 79.530 1.030 81.320 1.090 ;
        RECT 173.060 1.030 173.320 1.350 ;
        RECT 79.530 0.950 81.260 1.030 ;
        RECT 79.530 -4.800 80.090 0.950 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 102.190 1.600 102.510 1.660 ;
        RECT 195.570 1.600 195.890 1.660 ;
        RECT 102.190 1.460 195.890 1.600 ;
        RECT 102.190 1.400 102.510 1.460 ;
        RECT 195.570 1.400 195.890 1.460 ;
      LAYER met2 ;
        RECT 195.890 14.010 196.030 15.300 ;
        RECT 195.660 13.870 196.030 14.010 ;
        RECT 102.990 1.770 103.550 2.400 ;
        RECT 102.280 1.690 103.550 1.770 ;
        RECT 195.660 1.690 195.800 13.870 ;
        RECT 102.220 1.630 103.550 1.690 ;
        RECT 102.220 1.370 102.480 1.630 ;
        RECT 102.990 -4.800 103.550 1.630 ;
        RECT 195.600 1.370 195.860 1.690 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 128.870 4.660 129.190 4.720 ;
        RECT 217.650 4.660 217.970 4.720 ;
        RECT 128.870 4.520 217.970 4.660 ;
        RECT 128.870 4.460 129.190 4.520 ;
        RECT 217.650 4.460 217.970 4.520 ;
      LAYER met2 ;
        RECT 217.970 14.010 218.110 15.300 ;
        RECT 217.740 13.870 218.110 14.010 ;
        RECT 217.740 4.750 217.880 13.870 ;
        RECT 128.900 4.430 129.160 4.750 ;
        RECT 217.680 4.430 217.940 4.750 ;
        RECT 126.450 1.770 127.010 2.400 ;
        RECT 128.960 1.770 129.100 4.430 ;
        RECT 126.450 1.630 129.100 1.770 ;
        RECT 126.450 -4.800 127.010 1.630 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 58.490 5.680 58.810 5.740 ;
        RECT 123.810 5.680 124.130 5.740 ;
        RECT 58.490 5.540 124.130 5.680 ;
        RECT 58.490 5.480 58.810 5.540 ;
        RECT 123.810 5.480 124.130 5.540 ;
      LAYER met2 ;
        RECT 124.130 14.010 124.270 15.300 ;
        RECT 123.900 13.870 124.270 14.010 ;
        RECT 123.900 5.770 124.040 13.870 ;
        RECT 58.520 5.450 58.780 5.770 ;
        RECT 123.840 5.450 124.100 5.770 ;
        RECT 58.580 4.605 58.720 5.450 ;
        RECT 26.310 4.235 26.590 4.605 ;
        RECT 58.510 4.235 58.790 4.605 ;
        RECT 26.380 2.400 26.520 4.235 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER met3 ;
        RECT 26.285 4.570 26.615 4.585 ;
        RECT 58.485 4.570 58.815 4.585 ;
        RECT 26.285 4.270 58.815 4.570 ;
        RECT 26.285 4.255 26.615 4.270 ;
        RECT 58.485 4.255 58.815 4.270 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 54.810 6.360 55.130 6.420 ;
        RECT 129.330 6.360 129.650 6.420 ;
        RECT 54.810 6.220 129.650 6.360 ;
        RECT 54.810 6.160 55.130 6.220 ;
        RECT 129.330 6.160 129.650 6.220 ;
      LAYER met2 ;
        RECT 129.650 14.010 129.790 15.300 ;
        RECT 129.420 13.870 129.790 14.010 ;
        RECT 129.420 6.450 129.560 13.870 ;
        RECT 54.840 6.130 55.100 6.450 ;
        RECT 129.360 6.130 129.620 6.450 ;
        RECT 54.900 5.285 55.040 6.130 ;
        RECT 32.290 4.915 32.570 5.285 ;
        RECT 54.830 4.915 55.110 5.285 ;
        RECT 32.360 2.400 32.500 4.915 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER met3 ;
        RECT 32.265 5.250 32.595 5.265 ;
        RECT 54.805 5.250 55.135 5.265 ;
        RECT 32.265 4.950 55.135 5.250 ;
        RECT 32.265 4.935 32.595 4.950 ;
        RECT 54.805 4.935 55.135 4.950 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 71.080 3390.270 161.080 3396.070 ;
      LAYER pwell ;
        RECT 71.080 3385.220 161.080 3390.020 ;
      LAYER nwell ;
        RECT 93.530 3376.320 96.930 3377.920 ;
        RECT 93.530 3376.315 96.210 3376.320 ;
      LAYER pwell ;
        RECT 94.210 3376.020 96.015 3376.025 ;
        RECT 94.210 3375.795 96.930 3376.020 ;
        RECT 93.725 3375.120 96.930 3375.795 ;
        RECT 93.725 3375.115 96.015 3375.120 ;
        RECT 93.870 3374.925 94.040 3375.115 ;
        RECT 101.080 3370.270 161.080 3375.070 ;
      LAYER nwell ;
        RECT 101.080 3364.220 161.080 3370.020 ;
        RECT 68.180 3354.440 85.930 3356.140 ;
        RECT 112.580 3355.870 159.380 3359.670 ;
      LAYER pwell ;
        RECT 112.580 3355.470 114.880 3355.570 ;
        RECT 115.080 3355.470 125.780 3355.570 ;
        RECT 125.980 3355.470 130.480 3355.570 ;
        RECT 130.680 3355.470 141.380 3355.570 ;
        RECT 141.580 3355.470 146.080 3355.570 ;
        RECT 146.280 3355.470 156.980 3355.570 ;
        RECT 157.180 3355.470 159.380 3355.570 ;
        RECT 69.460 3353.990 70.805 3354.195 ;
        RECT 68.180 3353.965 69.030 3353.990 ;
        RECT 69.460 3353.965 72.430 3353.990 ;
        RECT 73.775 3353.965 74.695 3354.185 ;
        RECT 80.775 3354.085 81.695 3354.195 ;
        RECT 79.360 3353.990 81.695 3354.085 ;
        RECT 79.360 3353.965 83.930 3353.990 ;
        RECT 84.370 3353.965 85.715 3354.195 ;
        RECT 68.180 3353.290 85.715 3353.965 ;
        RECT 68.975 3353.285 70.805 3353.290 ;
        RECT 72.415 3353.285 81.695 3353.290 ;
        RECT 83.885 3353.285 85.715 3353.290 ;
        RECT 69.115 3353.095 69.285 3353.285 ;
        RECT 72.555 3353.095 72.725 3353.285 ;
        RECT 84.025 3353.095 84.195 3353.285 ;
        RECT 112.580 3352.770 159.380 3355.470 ;
      LAYER nwell ;
        RECT 68.230 3350.880 69.130 3350.940 ;
        RECT 68.230 3349.275 70.690 3350.880 ;
        RECT 80.530 3350.410 81.530 3350.440 ;
        RECT 68.230 3349.240 69.080 3349.275 ;
      LAYER pwell ;
        RECT 68.230 3348.985 69.180 3348.990 ;
        RECT 68.230 3348.090 70.485 3348.985 ;
      LAYER nwell ;
        RECT 76.940 3348.805 83.740 3350.410 ;
        RECT 80.530 3348.790 81.530 3348.805 ;
      LAYER pwell ;
        RECT 69.135 3348.075 70.485 3348.090 ;
        RECT 77.175 3348.290 80.345 3348.515 ;
        RECT 77.175 3348.285 81.730 3348.290 ;
        RECT 82.200 3348.285 83.545 3348.515 ;
        RECT 69.265 3347.885 69.435 3348.075 ;
        RECT 77.175 3347.605 83.545 3348.285 ;
      LAYER nwell ;
        RECT 119.580 3348.170 123.110 3349.770 ;
        RECT 120.430 3348.165 123.110 3348.170 ;
      LAYER pwell ;
        RECT 121.110 3347.645 122.915 3347.875 ;
        RECT 120.625 3347.640 122.915 3347.645 ;
        RECT 77.275 3347.415 77.445 3347.605 ;
        RECT 80.330 3347.590 81.730 3347.605 ;
        RECT 81.855 3347.415 82.025 3347.605 ;
        RECT 119.960 3346.965 122.915 3347.640 ;
        RECT 119.960 3346.960 120.630 3346.965 ;
        RECT 120.770 3346.775 120.940 3346.965 ;
        RECT 71.045 3345.425 71.215 3345.615 ;
        RECT 71.330 3345.425 72.830 3345.440 ;
        RECT 81.795 3345.425 81.965 3345.615 ;
        RECT 82.080 3345.425 84.080 3345.440 ;
        RECT 85.565 3345.425 85.735 3345.615 ;
        RECT 69.995 3344.745 85.875 3345.425 ;
        RECT 69.995 3344.625 75.160 3344.745 ;
        RECT 69.995 3344.515 73.745 3344.625 ;
        RECT 79.825 3344.525 80.745 3344.745 ;
        RECT 82.080 3344.740 85.390 3344.745 ;
        RECT 84.045 3344.515 85.390 3344.740 ;
        RECT 127.030 3344.670 158.230 3347.370 ;
        RECT 127.030 3344.570 129.230 3344.670 ;
        RECT 129.430 3344.570 140.130 3344.670 ;
        RECT 140.330 3344.570 144.830 3344.670 ;
        RECT 145.030 3344.570 155.730 3344.670 ;
        RECT 155.930 3344.570 158.230 3344.670 ;
        RECT 71.330 3344.490 72.830 3344.515 ;
      LAYER nwell ;
        RECT 71.530 3344.225 72.380 3344.240 ;
        RECT 82.280 3344.225 84.080 3344.240 ;
        RECT 69.790 3342.620 86.070 3344.225 ;
        RECT 71.530 3342.590 72.380 3342.620 ;
        RECT 82.280 3342.590 84.230 3342.620 ;
        RECT 127.030 3340.470 158.230 3344.270 ;
        RECT 70.780 3337.070 95.480 3337.120 ;
        RECT 70.580 3335.420 95.480 3337.070 ;
      LAYER pwell ;
        RECT 70.580 3334.220 95.480 3335.220 ;
      LAYER nwell ;
        RECT 138.030 3334.770 140.880 3336.370 ;
        RECT 138.030 3334.765 140.250 3334.770 ;
      LAYER pwell ;
        RECT 138.710 3334.470 140.055 3334.475 ;
        RECT 138.710 3334.245 140.880 3334.470 ;
        RECT 70.915 3334.075 71.085 3334.220 ;
        RECT 75.015 3334.075 75.185 3334.220 ;
        RECT 79.115 3334.075 79.285 3334.220 ;
        RECT 83.515 3334.075 83.685 3334.220 ;
        RECT 87.615 3334.075 87.785 3334.220 ;
        RECT 91.715 3334.075 91.885 3334.220 ;
        RECT 138.225 3333.570 140.880 3334.245 ;
        RECT 138.225 3333.565 140.055 3333.570 ;
        RECT 138.365 3333.375 138.535 3333.565 ;
      LAYER nwell ;
        RECT 71.730 3333.070 88.080 3333.120 ;
        RECT 70.580 3331.420 88.080 3333.070 ;
        RECT 143.730 3332.470 145.880 3332.520 ;
      LAYER pwell ;
        RECT 70.580 3330.220 88.080 3331.220 ;
        RECT 70.915 3330.075 71.085 3330.220 ;
        RECT 74.715 3330.075 74.885 3330.220 ;
        RECT 83.960 3330.075 84.130 3330.220 ;
        RECT 86.615 3330.075 86.785 3330.220 ;
      LAYER nwell ;
        RECT 115.580 3328.370 117.980 3330.970 ;
        RECT 119.330 3328.370 123.530 3330.970 ;
        RECT 124.830 3328.370 129.030 3330.970 ;
        RECT 130.330 3328.320 132.730 3330.920 ;
        RECT 143.730 3330.870 158.120 3332.470 ;
        RECT 145.780 3330.865 158.120 3330.870 ;
        RECT 148.380 3330.820 150.480 3330.865 ;
      LAYER pwell ;
        RECT 143.730 3330.575 146.080 3330.620 ;
        RECT 143.730 3330.370 148.215 3330.575 ;
        RECT 143.730 3330.345 150.630 3330.370 ;
        RECT 154.090 3330.345 155.000 3330.565 ;
        RECT 156.535 3330.345 157.885 3330.575 ;
        RECT 143.730 3329.665 157.885 3330.345 ;
        RECT 143.730 3329.620 146.080 3329.665 ;
        RECT 146.115 3329.475 146.285 3329.665 ;
        RECT 148.180 3329.620 150.630 3329.665 ;
        RECT 150.715 3329.475 150.885 3329.665 ;
      LAYER nwell ;
        RECT 142.730 3326.670 160.480 3328.270 ;
        RECT 143.580 3326.665 160.480 3326.670 ;
        RECT 146.680 3326.620 149.030 3326.665 ;
        RECT 158.980 3326.620 160.480 3326.665 ;
      LAYER pwell ;
        RECT 143.775 3326.370 146.385 3326.375 ;
        RECT 142.730 3326.170 146.385 3326.370 ;
        RECT 142.730 3326.145 149.230 3326.170 ;
        RECT 152.690 3326.145 153.600 3326.365 ;
        RECT 155.140 3326.145 158.825 3326.375 ;
        RECT 142.730 3325.465 158.825 3326.145 ;
        RECT 142.730 3325.120 143.830 3325.465 ;
        RECT 143.920 3325.275 144.090 3325.465 ;
        RECT 146.380 3325.420 149.230 3325.465 ;
        RECT 149.315 3325.275 149.485 3325.465 ;
        RECT 158.830 3325.420 160.480 3326.370 ;
      LAYER nwell ;
        RECT 68.180 3322.790 85.930 3324.490 ;
      LAYER pwell ;
        RECT 69.460 3322.340 70.805 3322.545 ;
        RECT 68.180 3322.315 69.030 3322.340 ;
        RECT 69.460 3322.315 72.430 3322.340 ;
        RECT 73.775 3322.315 74.695 3322.535 ;
        RECT 80.775 3322.435 81.695 3322.545 ;
        RECT 79.360 3322.340 81.695 3322.435 ;
        RECT 79.360 3322.315 83.930 3322.340 ;
        RECT 84.370 3322.315 85.715 3322.545 ;
        RECT 68.180 3321.640 85.715 3322.315 ;
        RECT 68.975 3321.635 70.805 3321.640 ;
        RECT 72.415 3321.635 81.695 3321.640 ;
        RECT 83.885 3321.635 85.715 3321.640 ;
        RECT 69.115 3321.445 69.285 3321.635 ;
        RECT 72.555 3321.445 72.725 3321.635 ;
        RECT 84.025 3321.445 84.195 3321.635 ;
        RECT 109.525 3321.185 110.205 3321.325 ;
        RECT 109.335 3321.015 110.205 3321.185 ;
        RECT 109.525 3320.840 110.205 3321.015 ;
        RECT 109.525 3319.495 110.435 3320.840 ;
      LAYER nwell ;
        RECT 68.230 3319.230 69.130 3319.290 ;
        RECT 68.230 3317.625 70.690 3319.230 ;
        RECT 80.530 3318.760 81.530 3318.790 ;
        RECT 68.230 3317.590 69.080 3317.625 ;
      LAYER pwell ;
        RECT 68.230 3317.335 69.180 3317.340 ;
        RECT 68.230 3316.440 70.485 3317.335 ;
      LAYER nwell ;
        RECT 76.940 3317.155 83.740 3318.760 ;
      LAYER pwell ;
        RECT 109.530 3318.015 110.430 3319.495 ;
      LAYER nwell ;
        RECT 110.725 3319.370 112.330 3321.520 ;
        RECT 110.680 3318.220 112.330 3319.370 ;
        RECT 115.930 3319.120 119.230 3323.920 ;
      LAYER pwell ;
        RECT 120.730 3320.970 124.030 3323.770 ;
        RECT 125.280 3320.970 128.580 3323.770 ;
      LAYER nwell ;
        RECT 129.780 3319.070 133.080 3323.870 ;
        RECT 143.730 3320.770 145.880 3320.820 ;
        RECT 143.730 3319.170 158.120 3320.770 ;
        RECT 145.780 3319.165 158.120 3319.170 ;
        RECT 148.380 3319.120 150.480 3319.165 ;
      LAYER pwell ;
        RECT 109.525 3317.885 110.435 3318.015 ;
        RECT 109.335 3317.715 110.435 3317.885 ;
      LAYER nwell ;
        RECT 80.530 3317.140 81.530 3317.155 ;
      LAYER pwell ;
        RECT 69.135 3316.425 70.485 3316.440 ;
        RECT 77.175 3316.640 80.345 3316.865 ;
        RECT 77.175 3316.635 81.730 3316.640 ;
        RECT 82.200 3316.635 83.545 3316.865 ;
        RECT 109.525 3316.665 110.435 3317.715 ;
        RECT 69.265 3316.235 69.435 3316.425 ;
        RECT 77.175 3315.955 83.545 3316.635 ;
      LAYER nwell ;
        RECT 110.725 3316.460 112.330 3318.220 ;
      LAYER pwell ;
        RECT 143.730 3318.875 146.080 3318.920 ;
        RECT 143.730 3318.670 148.215 3318.875 ;
        RECT 143.730 3318.645 150.630 3318.670 ;
        RECT 154.090 3318.645 155.000 3318.865 ;
        RECT 156.535 3318.645 157.885 3318.875 ;
        RECT 143.730 3317.965 157.885 3318.645 ;
        RECT 143.730 3317.920 146.080 3317.965 ;
        RECT 146.115 3317.775 146.285 3317.965 ;
        RECT 148.180 3317.920 150.630 3317.965 ;
        RECT 150.715 3317.775 150.885 3317.965 ;
        RECT 77.275 3315.765 77.445 3315.955 ;
        RECT 80.330 3315.940 81.730 3315.955 ;
        RECT 81.855 3315.765 82.025 3315.955 ;
        RECT 71.045 3313.775 71.215 3313.965 ;
        RECT 71.330 3313.775 72.830 3313.790 ;
        RECT 81.795 3313.775 81.965 3313.965 ;
        RECT 82.080 3313.775 84.080 3313.790 ;
        RECT 85.565 3313.775 85.735 3313.965 ;
        RECT 69.995 3313.095 85.875 3313.775 ;
        RECT 69.995 3312.975 75.160 3313.095 ;
        RECT 69.995 3312.865 73.745 3312.975 ;
        RECT 79.825 3312.875 80.745 3313.095 ;
        RECT 82.080 3313.090 85.390 3313.095 ;
        RECT 84.045 3312.865 85.390 3313.090 ;
        RECT 118.180 3312.970 132.560 3314.980 ;
      LAYER nwell ;
        RECT 142.730 3314.970 160.480 3316.570 ;
        RECT 143.580 3314.965 160.480 3314.970 ;
        RECT 146.680 3314.920 149.030 3314.965 ;
        RECT 158.980 3314.920 160.480 3314.965 ;
      LAYER pwell ;
        RECT 143.775 3314.670 146.385 3314.675 ;
        RECT 142.730 3314.470 146.385 3314.670 ;
        RECT 142.730 3314.445 149.230 3314.470 ;
        RECT 152.690 3314.445 153.600 3314.665 ;
        RECT 155.140 3314.445 158.825 3314.675 ;
        RECT 142.730 3313.765 158.825 3314.445 ;
        RECT 142.730 3313.420 143.830 3313.765 ;
        RECT 143.920 3313.575 144.090 3313.765 ;
        RECT 146.380 3313.720 149.230 3313.765 ;
        RECT 149.315 3313.575 149.485 3313.765 ;
        RECT 158.830 3313.720 160.480 3314.670 ;
        RECT 71.330 3312.840 72.830 3312.865 ;
      LAYER nwell ;
        RECT 71.530 3312.575 72.380 3312.590 ;
        RECT 82.280 3312.575 84.080 3312.590 ;
        RECT 69.790 3310.970 86.070 3312.575 ;
        RECT 71.530 3310.940 72.380 3310.970 ;
        RECT 82.280 3310.940 84.230 3310.970 ;
      LAYER li1 ;
        RECT 71.280 3396.570 171.280 3396.970 ;
        RECT 71.280 3395.220 71.680 3396.570 ;
        RECT 71.980 3390.670 72.380 3396.570 ;
        RECT 73.180 3389.820 74.380 3390.470 ;
        RECT 71.280 3385.570 71.680 3386.070 ;
        RECT 71.980 3384.720 72.380 3389.620 ;
        RECT 76.030 3389.270 76.430 3395.670 ;
        RECT 80.080 3390.670 80.480 3396.570 ;
        RECT 80.780 3395.670 81.180 3396.570 ;
        RECT 81.480 3395.670 81.880 3396.570 ;
        RECT 86.230 3395.670 86.630 3396.570 ;
        RECT 86.930 3395.670 87.330 3396.570 ;
        RECT 80.780 3395.220 81.880 3395.670 ;
        RECT 81.480 3390.670 81.880 3395.220 ;
        RECT 76.880 3389.820 78.080 3390.470 ;
        RECT 83.030 3390.370 84.230 3390.470 ;
        RECT 78.880 3389.870 84.230 3390.370 ;
        RECT 78.880 3389.270 79.380 3389.870 ;
        RECT 83.030 3389.820 84.230 3389.870 ;
        RECT 85.530 3390.420 85.930 3395.670 ;
        RECT 86.230 3395.220 87.330 3395.670 ;
        RECT 86.930 3390.670 87.330 3395.220 ;
        RECT 87.880 3390.420 89.080 3390.470 ;
        RECT 85.530 3389.920 89.080 3390.420 ;
        RECT 76.030 3388.770 79.380 3389.270 ;
        RECT 76.030 3385.620 76.430 3388.770 ;
        RECT 80.080 3384.720 80.480 3389.620 ;
        RECT 80.780 3385.570 81.180 3386.070 ;
        RECT 81.480 3384.720 81.880 3389.620 ;
        RECT 85.530 3385.620 85.930 3389.920 ;
        RECT 87.880 3389.820 89.080 3389.920 ;
        RECT 86.230 3385.570 86.630 3386.070 ;
        RECT 86.930 3384.720 87.330 3389.620 ;
        RECT 90.980 3385.620 91.380 3395.670 ;
        RECT 91.680 3395.220 92.080 3396.570 ;
        RECT 92.380 3390.670 92.780 3396.570 ;
        RECT 93.580 3389.820 94.780 3390.470 ;
        RECT 91.680 3385.570 92.080 3386.070 ;
        RECT 92.380 3384.720 92.780 3389.620 ;
        RECT 96.430 3385.620 96.830 3395.670 ;
        RECT 100.480 3390.670 100.880 3396.570 ;
        RECT 101.280 3395.220 101.680 3396.570 ;
        RECT 101.980 3390.670 102.380 3396.570 ;
        RECT 97.280 3389.820 98.480 3390.470 ;
        RECT 103.180 3389.820 104.380 3390.470 ;
        RECT 100.480 3384.720 100.880 3389.620 ;
        RECT 101.280 3385.570 101.680 3386.070 ;
        RECT 101.980 3384.720 102.380 3389.620 ;
        RECT 106.030 3389.270 106.430 3395.670 ;
        RECT 110.080 3390.670 110.480 3396.570 ;
        RECT 110.780 3395.670 111.180 3396.570 ;
        RECT 111.480 3395.670 111.880 3396.570 ;
        RECT 116.230 3395.670 116.630 3396.570 ;
        RECT 116.930 3395.670 117.330 3396.570 ;
        RECT 110.780 3395.220 111.880 3395.670 ;
        RECT 111.480 3390.670 111.880 3395.220 ;
        RECT 106.880 3389.820 108.080 3390.470 ;
        RECT 113.030 3390.370 114.230 3390.470 ;
        RECT 108.880 3389.870 114.230 3390.370 ;
        RECT 108.880 3389.270 109.380 3389.870 ;
        RECT 113.030 3389.820 114.230 3389.870 ;
        RECT 115.530 3390.420 115.930 3395.670 ;
        RECT 116.230 3395.220 117.330 3395.670 ;
        RECT 116.930 3390.670 117.330 3395.220 ;
        RECT 117.880 3390.420 119.080 3390.470 ;
        RECT 115.530 3389.920 119.080 3390.420 ;
        RECT 106.030 3388.770 109.380 3389.270 ;
        RECT 106.030 3385.620 106.430 3388.770 ;
        RECT 110.080 3384.720 110.480 3389.620 ;
        RECT 110.780 3385.570 111.180 3386.070 ;
        RECT 111.480 3384.720 111.880 3389.620 ;
        RECT 115.530 3385.620 115.930 3389.920 ;
        RECT 117.880 3389.820 119.080 3389.920 ;
        RECT 116.230 3385.570 116.630 3386.070 ;
        RECT 116.930 3384.720 117.330 3389.620 ;
        RECT 120.980 3385.620 121.380 3395.670 ;
        RECT 121.680 3395.220 122.080 3396.570 ;
        RECT 122.380 3390.670 122.780 3396.570 ;
        RECT 123.580 3389.820 124.780 3390.470 ;
        RECT 121.680 3385.570 122.080 3386.070 ;
        RECT 122.380 3384.720 122.780 3389.620 ;
        RECT 126.430 3385.620 126.830 3395.670 ;
        RECT 130.480 3390.670 130.880 3396.570 ;
        RECT 131.280 3395.220 131.680 3396.570 ;
        RECT 131.980 3390.670 132.380 3396.570 ;
        RECT 127.280 3389.820 128.480 3390.470 ;
        RECT 133.180 3389.820 134.380 3390.470 ;
        RECT 130.480 3384.720 130.880 3389.620 ;
        RECT 131.280 3385.570 131.680 3386.070 ;
        RECT 131.980 3384.720 132.380 3389.620 ;
        RECT 136.030 3389.270 136.430 3395.670 ;
        RECT 140.080 3390.670 140.480 3396.570 ;
        RECT 140.780 3395.670 141.180 3396.570 ;
        RECT 141.480 3395.670 141.880 3396.570 ;
        RECT 146.230 3395.670 146.630 3396.570 ;
        RECT 146.930 3395.670 147.330 3396.570 ;
        RECT 140.780 3395.220 141.880 3395.670 ;
        RECT 141.480 3390.670 141.880 3395.220 ;
        RECT 136.880 3389.820 138.080 3390.470 ;
        RECT 143.030 3390.370 144.230 3390.470 ;
        RECT 138.880 3389.870 144.230 3390.370 ;
        RECT 138.880 3389.270 139.380 3389.870 ;
        RECT 143.030 3389.820 144.230 3389.870 ;
        RECT 145.530 3390.420 145.930 3395.670 ;
        RECT 146.230 3395.220 147.330 3395.670 ;
        RECT 146.930 3390.670 147.330 3395.220 ;
        RECT 147.880 3390.420 149.080 3390.470 ;
        RECT 145.530 3389.920 149.080 3390.420 ;
        RECT 136.030 3388.770 139.380 3389.270 ;
        RECT 136.030 3385.620 136.430 3388.770 ;
        RECT 140.080 3384.720 140.480 3389.620 ;
        RECT 140.780 3385.570 141.180 3386.070 ;
        RECT 141.480 3384.720 141.880 3389.620 ;
        RECT 145.530 3385.620 145.930 3389.920 ;
        RECT 147.880 3389.820 149.080 3389.920 ;
        RECT 146.230 3385.570 146.630 3386.070 ;
        RECT 146.930 3384.720 147.330 3389.620 ;
        RECT 150.980 3385.620 151.380 3395.670 ;
        RECT 151.680 3395.220 152.080 3396.570 ;
        RECT 152.380 3390.670 152.780 3396.570 ;
        RECT 153.580 3389.820 154.780 3390.470 ;
        RECT 151.680 3385.570 152.080 3386.070 ;
        RECT 152.380 3384.720 152.780 3389.620 ;
        RECT 156.430 3385.620 156.830 3395.670 ;
        RECT 160.480 3390.670 160.880 3396.570 ;
        RECT 157.280 3389.820 158.480 3390.470 ;
        RECT 160.480 3384.720 160.880 3389.620 ;
        RECT 71.980 3384.320 160.880 3384.720 ;
        RECT 102.030 3381.270 102.530 3384.320 ;
        RECT 102.930 3381.270 103.380 3381.320 ;
        RECT 102.030 3381.220 103.380 3381.270 ;
        RECT 102.030 3380.900 105.195 3381.220 ;
        RECT 102.030 3380.870 103.380 3380.900 ;
        RECT 102.030 3379.820 102.530 3380.870 ;
        RECT 102.930 3380.820 103.380 3380.870 ;
        RECT 102.030 3379.750 103.280 3379.820 ;
        RECT 102.030 3379.670 103.380 3379.750 ;
        RECT 109.180 3379.670 109.350 3379.750 ;
        RECT 102.030 3379.350 105.195 3379.670 ;
        RECT 107.365 3379.350 109.350 3379.670 ;
        RECT 102.030 3379.270 103.380 3379.350 ;
        RECT 109.180 3379.270 109.350 3379.350 ;
        RECT 102.030 3379.220 103.280 3379.270 ;
        RECT 93.720 3377.645 96.020 3377.815 ;
        RECT 93.805 3377.075 94.065 3377.475 ;
        RECT 94.235 3377.245 95.170 3377.645 ;
        RECT 95.340 3377.135 95.935 3377.475 ;
        RECT 64.180 3376.070 73.030 3377.070 ;
        RECT 87.430 3376.070 88.430 3377.070 ;
        RECT 93.805 3376.905 95.170 3377.075 ;
        RECT 92.530 3376.670 93.430 3376.770 ;
        RECT 93.805 3376.670 94.265 3376.735 ;
        RECT 92.530 3376.370 94.265 3376.670 ;
        RECT 92.530 3376.270 93.430 3376.370 ;
        RECT 87.630 3363.470 88.180 3376.070 ;
        RECT 93.805 3376.005 94.265 3376.370 ;
        RECT 94.435 3375.835 95.170 3376.905 ;
        RECT 93.805 3375.665 95.170 3375.835 ;
        RECT 95.340 3375.815 95.515 3377.135 ;
        RECT 95.695 3376.670 95.935 3376.965 ;
        RECT 96.280 3376.870 96.680 3377.370 ;
        RECT 95.695 3376.170 96.130 3376.670 ;
        RECT 95.695 3375.985 95.935 3376.170 ;
        RECT 93.805 3375.265 94.065 3375.665 ;
        RECT 94.235 3375.095 95.170 3375.495 ;
        RECT 95.340 3375.265 95.935 3375.815 ;
        RECT 96.280 3375.370 96.680 3375.870 ;
        RECT 93.720 3374.925 96.020 3375.095 ;
        RECT 97.330 3363.720 97.830 3376.670 ;
        RECT 102.030 3375.970 102.530 3379.220 ;
        RECT 159.680 3375.970 160.180 3384.320 ;
        RECT 101.280 3375.570 160.180 3375.970 ;
        RECT 101.280 3370.670 101.680 3375.570 ;
        RECT 103.680 3369.820 104.880 3370.470 ;
        RECT 101.280 3363.720 101.680 3369.620 ;
        RECT 105.330 3364.620 105.730 3374.670 ;
        RECT 109.380 3370.670 109.780 3375.570 ;
        RECT 110.080 3374.220 110.480 3374.720 ;
        RECT 107.380 3369.820 108.580 3370.470 ;
        RECT 109.380 3363.720 109.780 3369.620 ;
        RECT 110.080 3363.720 110.480 3365.070 ;
        RECT 110.780 3364.620 111.180 3374.670 ;
        RECT 114.830 3370.670 115.230 3375.570 ;
        RECT 115.530 3374.220 115.930 3374.720 ;
        RECT 113.080 3370.370 114.280 3370.470 ;
        RECT 116.230 3370.370 116.630 3374.670 ;
        RECT 120.280 3370.670 120.680 3375.570 ;
        RECT 120.980 3374.220 121.380 3374.720 ;
        RECT 121.680 3370.670 122.080 3375.570 ;
        RECT 125.730 3371.520 126.130 3374.670 ;
        RECT 122.780 3371.020 126.130 3371.520 ;
        RECT 113.080 3369.870 116.630 3370.370 ;
        RECT 113.080 3369.820 114.280 3369.870 ;
        RECT 114.830 3365.070 115.230 3369.620 ;
        RECT 114.830 3364.620 115.930 3365.070 ;
        RECT 116.230 3364.620 116.630 3369.870 ;
        RECT 117.930 3370.420 119.130 3370.470 ;
        RECT 122.780 3370.420 123.280 3371.020 ;
        RECT 117.930 3369.920 123.280 3370.420 ;
        RECT 117.930 3369.820 119.130 3369.920 ;
        RECT 124.080 3369.820 125.280 3370.470 ;
        RECT 120.280 3365.070 120.680 3369.620 ;
        RECT 120.280 3364.620 121.380 3365.070 ;
        RECT 114.830 3363.720 115.230 3364.620 ;
        RECT 115.530 3363.720 115.930 3364.620 ;
        RECT 120.280 3363.720 120.680 3364.620 ;
        RECT 120.980 3363.720 121.380 3364.620 ;
        RECT 121.680 3363.720 122.080 3369.620 ;
        RECT 125.730 3364.620 126.130 3371.020 ;
        RECT 129.780 3370.670 130.180 3375.570 ;
        RECT 130.480 3374.220 130.880 3374.720 ;
        RECT 131.280 3370.670 131.680 3375.570 ;
        RECT 127.780 3369.820 128.980 3370.470 ;
        RECT 133.680 3369.820 134.880 3370.470 ;
        RECT 129.780 3363.720 130.180 3369.620 ;
        RECT 130.480 3363.720 130.880 3365.070 ;
        RECT 131.280 3363.720 131.680 3369.620 ;
        RECT 135.330 3364.620 135.730 3374.670 ;
        RECT 139.380 3370.670 139.780 3375.570 ;
        RECT 140.080 3374.220 140.480 3374.720 ;
        RECT 137.380 3369.820 138.580 3370.470 ;
        RECT 139.380 3363.720 139.780 3369.620 ;
        RECT 140.080 3363.720 140.480 3365.070 ;
        RECT 140.780 3364.620 141.180 3374.670 ;
        RECT 144.830 3370.670 145.230 3375.570 ;
        RECT 145.530 3374.220 145.930 3374.720 ;
        RECT 143.080 3370.370 144.280 3370.470 ;
        RECT 146.230 3370.370 146.630 3374.670 ;
        RECT 150.280 3370.670 150.680 3375.570 ;
        RECT 150.980 3374.220 151.380 3374.720 ;
        RECT 151.680 3370.670 152.080 3375.570 ;
        RECT 155.730 3371.520 156.130 3374.670 ;
        RECT 152.780 3371.020 156.130 3371.520 ;
        RECT 143.080 3369.870 146.630 3370.370 ;
        RECT 143.080 3369.820 144.280 3369.870 ;
        RECT 144.830 3365.070 145.230 3369.620 ;
        RECT 144.830 3364.620 145.930 3365.070 ;
        RECT 146.230 3364.620 146.630 3369.870 ;
        RECT 147.930 3370.420 149.130 3370.470 ;
        RECT 152.780 3370.420 153.280 3371.020 ;
        RECT 147.930 3369.920 153.280 3370.420 ;
        RECT 147.930 3369.820 149.130 3369.920 ;
        RECT 154.080 3369.820 155.280 3370.470 ;
        RECT 150.280 3365.070 150.680 3369.620 ;
        RECT 150.280 3364.620 151.380 3365.070 ;
        RECT 144.830 3363.720 145.230 3364.620 ;
        RECT 145.530 3363.720 145.930 3364.620 ;
        RECT 150.280 3363.720 150.680 3364.620 ;
        RECT 150.980 3363.720 151.380 3364.620 ;
        RECT 151.680 3363.720 152.080 3369.620 ;
        RECT 155.730 3364.620 156.130 3371.020 ;
        RECT 159.780 3370.670 160.180 3375.570 ;
        RECT 160.480 3374.220 160.880 3374.720 ;
        RECT 157.780 3369.820 158.980 3370.470 ;
        RECT 159.780 3363.720 160.180 3369.620 ;
        RECT 160.480 3363.720 160.880 3365.070 ;
        RECT 170.280 3363.720 171.280 3396.570 ;
        RECT 97.330 3363.320 171.280 3363.720 ;
        RECT 97.330 3363.220 101.680 3363.320 ;
        RECT 112.780 3360.170 159.180 3360.570 ;
        RECT 112.780 3358.820 113.180 3360.170 ;
        RECT 113.480 3356.270 113.880 3360.170 ;
        RECT 85.630 3355.985 88.180 3355.990 ;
        RECT 68.970 3355.815 70.810 3355.985 ;
        RECT 72.410 3355.815 82.070 3355.985 ;
        RECT 83.880 3355.815 88.180 3355.985 ;
        RECT 69.145 3354.885 69.315 3355.645 ;
        RECT 69.530 3355.055 69.860 3355.815 ;
        RECT 69.145 3354.715 69.860 3354.885 ;
        RECT 70.030 3354.740 70.285 3355.645 ;
        RECT 68.080 3354.190 69.430 3354.540 ;
        RECT 69.690 3354.505 69.860 3354.715 ;
        RECT 69.055 3354.165 69.410 3354.190 ;
        RECT 69.690 3354.175 69.945 3354.505 ;
        RECT 70.115 3354.490 70.285 3354.740 ;
        RECT 70.460 3354.665 70.720 3355.815 ;
        RECT 71.430 3355.040 71.830 3355.540 ;
        RECT 72.585 3355.145 72.755 3355.645 ;
        RECT 72.925 3355.315 73.255 3355.815 ;
        RECT 72.585 3354.975 73.250 3355.145 ;
        RECT 72.500 3354.490 72.850 3354.805 ;
        RECT 70.115 3354.290 72.850 3354.490 ;
        RECT 69.690 3353.985 69.860 3354.175 ;
        RECT 70.115 3354.010 70.285 3354.290 ;
        RECT 72.500 3354.155 72.850 3354.290 ;
        RECT 68.380 3353.440 68.780 3353.940 ;
        RECT 69.145 3353.815 69.860 3353.985 ;
        RECT 69.145 3353.435 69.315 3353.815 ;
        RECT 69.530 3353.265 69.860 3353.645 ;
        RECT 70.030 3353.435 70.285 3354.010 ;
        RECT 70.460 3353.440 70.720 3354.105 ;
        RECT 73.020 3353.985 73.250 3354.975 ;
        RECT 72.585 3353.815 73.250 3353.985 ;
        RECT 72.585 3353.525 72.755 3353.815 ;
        RECT 70.460 3353.265 72.430 3353.440 ;
        RECT 72.925 3353.265 73.255 3353.645 ;
        RECT 73.425 3353.525 73.650 3355.645 ;
        RECT 73.865 3355.315 74.195 3355.815 ;
        RECT 74.365 3355.145 74.535 3355.645 ;
        RECT 74.770 3355.430 75.600 3355.600 ;
        RECT 75.840 3355.435 76.220 3355.815 ;
        RECT 73.840 3354.975 74.535 3355.145 ;
        RECT 73.840 3354.005 74.010 3354.975 ;
        RECT 74.180 3354.185 74.590 3354.805 ;
        RECT 74.760 3354.755 75.260 3355.135 ;
        RECT 73.840 3353.815 74.535 3354.005 ;
        RECT 74.760 3353.885 74.980 3354.755 ;
        RECT 75.430 3354.585 75.600 3355.430 ;
        RECT 76.400 3355.265 76.570 3355.555 ;
        RECT 76.740 3355.435 77.070 3355.815 ;
        RECT 77.540 3355.345 78.170 3355.595 ;
        RECT 78.350 3355.435 78.770 3355.815 ;
        RECT 78.000 3355.265 78.170 3355.345 ;
        RECT 78.970 3355.265 79.210 3355.555 ;
        RECT 75.770 3355.015 77.140 3355.265 ;
        RECT 75.770 3354.755 76.020 3355.015 ;
        RECT 76.530 3354.585 76.780 3354.745 ;
        RECT 75.430 3354.415 76.780 3354.585 ;
        RECT 75.430 3354.375 75.850 3354.415 ;
        RECT 75.160 3353.825 75.510 3354.195 ;
        RECT 73.865 3353.265 74.195 3353.645 ;
        RECT 74.365 3353.485 74.535 3353.815 ;
        RECT 75.680 3353.645 75.850 3354.375 ;
        RECT 76.950 3354.245 77.140 3355.015 ;
        RECT 76.020 3353.915 76.430 3354.245 ;
        RECT 76.720 3353.905 77.140 3354.245 ;
        RECT 77.310 3354.835 77.830 3355.145 ;
        RECT 78.000 3355.095 79.210 3355.265 ;
        RECT 79.440 3355.125 79.770 3355.815 ;
        RECT 77.310 3354.075 77.480 3354.835 ;
        RECT 77.650 3354.245 77.830 3354.655 ;
        RECT 78.000 3354.585 78.170 3355.095 ;
        RECT 79.940 3354.945 80.110 3355.555 ;
        RECT 80.380 3355.095 80.710 3355.605 ;
        RECT 79.940 3354.925 80.260 3354.945 ;
        RECT 78.340 3354.755 80.260 3354.925 ;
        RECT 78.000 3354.415 79.900 3354.585 ;
        RECT 78.230 3354.075 78.560 3354.195 ;
        RECT 77.310 3353.905 78.560 3354.075 ;
        RECT 74.835 3353.445 75.850 3353.645 ;
        RECT 76.020 3353.265 76.430 3353.705 ;
        RECT 76.720 3353.475 76.970 3353.905 ;
        RECT 77.170 3353.265 77.490 3353.725 ;
        RECT 78.730 3353.655 78.900 3354.415 ;
        RECT 79.570 3354.355 79.900 3354.415 ;
        RECT 79.090 3354.185 79.420 3354.245 ;
        RECT 79.090 3353.915 79.750 3354.185 ;
        RECT 80.070 3353.860 80.260 3354.755 ;
        RECT 78.050 3353.485 78.900 3353.655 ;
        RECT 79.100 3353.265 79.760 3353.745 ;
        RECT 79.940 3353.530 80.260 3353.860 ;
        RECT 80.460 3354.505 80.710 3355.095 ;
        RECT 80.890 3355.015 81.175 3355.815 ;
        RECT 81.355 3354.835 81.610 3355.505 ;
        RECT 81.430 3354.540 81.610 3354.835 ;
        RECT 84.055 3354.885 84.225 3355.645 ;
        RECT 84.440 3355.055 84.770 3355.815 ;
        RECT 84.055 3354.715 84.770 3354.885 ;
        RECT 84.940 3354.740 85.195 3355.645 ;
        RECT 81.430 3354.535 83.980 3354.540 ;
        RECT 80.460 3354.175 81.260 3354.505 ;
        RECT 80.460 3353.525 80.710 3354.175 ;
        RECT 81.430 3354.165 84.320 3354.535 ;
        RECT 84.600 3354.505 84.770 3354.715 ;
        RECT 84.600 3354.175 84.855 3354.505 ;
        RECT 81.430 3354.140 83.980 3354.165 ;
        RECT 81.430 3353.975 81.610 3354.140 ;
        RECT 84.600 3353.985 84.770 3354.175 ;
        RECT 85.025 3354.010 85.195 3354.740 ;
        RECT 85.370 3355.640 88.180 3355.815 ;
        RECT 85.370 3354.665 85.630 3355.640 ;
        RECT 87.830 3355.190 88.180 3355.640 ;
        RECT 114.130 3355.470 114.580 3355.920 ;
        RECT 80.890 3353.265 81.175 3353.725 ;
        RECT 81.355 3353.445 81.610 3353.975 ;
        RECT 84.055 3353.815 84.770 3353.985 ;
        RECT 84.055 3353.435 84.225 3353.815 ;
        RECT 82.030 3353.265 83.880 3353.390 ;
        RECT 84.440 3353.265 84.770 3353.645 ;
        RECT 84.940 3353.435 85.195 3354.010 ;
        RECT 85.370 3353.265 85.630 3354.105 ;
        RECT 68.970 3353.095 85.720 3353.265 ;
        RECT 70.680 3352.940 72.430 3353.095 ;
        RECT 82.030 3352.940 83.880 3353.095 ;
        RECT 112.780 3352.270 113.180 3353.620 ;
        RECT 113.480 3352.270 113.880 3355.170 ;
        RECT 115.080 3353.170 115.480 3359.270 ;
        RECT 116.680 3356.270 117.080 3360.170 ;
        RECT 117.480 3359.220 117.880 3360.170 ;
        RECT 118.180 3359.220 118.580 3359.270 ;
        RECT 117.480 3358.720 118.580 3359.220 ;
        RECT 118.180 3356.270 118.580 3358.720 ;
        RECT 119.780 3355.970 120.180 3359.270 ;
        RECT 120.580 3359.220 120.980 3360.170 ;
        RECT 121.280 3359.220 121.680 3359.270 ;
        RECT 120.580 3358.720 121.680 3359.220 ;
        RECT 121.280 3356.270 121.680 3358.720 ;
        RECT 115.730 3355.470 116.180 3355.920 ;
        RECT 118.580 3355.470 119.530 3355.970 ;
        RECT 119.780 3355.470 122.630 3355.970 ;
        RECT 116.680 3352.270 117.080 3355.170 ;
        RECT 118.180 3353.620 118.580 3355.170 ;
        RECT 117.480 3353.170 118.580 3353.620 ;
        RECT 119.780 3353.170 120.180 3355.470 ;
        RECT 121.280 3353.620 121.680 3355.170 ;
        RECT 120.580 3353.170 121.680 3353.620 ;
        RECT 122.880 3353.170 123.280 3359.270 ;
        RECT 123.680 3358.820 124.080 3360.170 ;
        RECT 124.380 3356.270 124.780 3360.170 ;
        RECT 125.030 3355.470 125.480 3355.920 ;
        RECT 117.480 3353.120 117.880 3353.170 ;
        RECT 118.180 3352.270 118.580 3353.170 ;
        RECT 120.580 3353.120 120.980 3353.170 ;
        RECT 121.280 3352.270 121.680 3353.170 ;
        RECT 123.680 3352.270 124.080 3353.620 ;
        RECT 124.380 3352.270 124.780 3355.170 ;
        RECT 125.980 3353.170 126.380 3359.270 ;
        RECT 127.580 3356.270 127.980 3360.170 ;
        RECT 128.380 3358.820 128.780 3360.170 ;
        RECT 129.080 3356.270 129.480 3360.170 ;
        RECT 126.630 3355.470 127.080 3355.920 ;
        RECT 129.730 3355.470 130.180 3355.920 ;
        RECT 127.580 3352.270 127.980 3355.170 ;
        RECT 128.380 3352.270 128.780 3353.620 ;
        RECT 129.080 3352.270 129.480 3355.170 ;
        RECT 130.680 3353.170 131.080 3359.270 ;
        RECT 132.280 3356.270 132.680 3360.170 ;
        RECT 133.080 3359.220 133.480 3360.170 ;
        RECT 133.780 3359.220 134.180 3359.270 ;
        RECT 133.080 3358.720 134.180 3359.220 ;
        RECT 133.780 3356.270 134.180 3358.720 ;
        RECT 135.380 3355.970 135.780 3359.270 ;
        RECT 136.180 3359.220 136.580 3360.170 ;
        RECT 136.880 3359.220 137.280 3359.270 ;
        RECT 136.180 3358.720 137.280 3359.220 ;
        RECT 136.880 3356.270 137.280 3358.720 ;
        RECT 131.330 3355.470 131.780 3355.920 ;
        RECT 134.180 3355.470 135.130 3355.970 ;
        RECT 135.380 3355.470 138.230 3355.970 ;
        RECT 132.280 3352.270 132.680 3355.170 ;
        RECT 133.780 3353.620 134.180 3355.170 ;
        RECT 133.080 3353.170 134.180 3353.620 ;
        RECT 135.380 3353.170 135.780 3355.470 ;
        RECT 136.880 3353.620 137.280 3355.170 ;
        RECT 136.180 3353.170 137.280 3353.620 ;
        RECT 138.480 3353.170 138.880 3359.270 ;
        RECT 139.280 3358.820 139.680 3360.170 ;
        RECT 139.980 3356.270 140.380 3360.170 ;
        RECT 140.630 3355.470 141.080 3355.920 ;
        RECT 133.080 3353.120 133.480 3353.170 ;
        RECT 133.780 3352.270 134.180 3353.170 ;
        RECT 136.180 3353.120 136.580 3353.170 ;
        RECT 136.880 3352.270 137.280 3353.170 ;
        RECT 139.280 3352.270 139.680 3353.620 ;
        RECT 139.980 3352.270 140.380 3355.170 ;
        RECT 141.580 3353.170 141.980 3359.270 ;
        RECT 143.180 3356.270 143.580 3360.170 ;
        RECT 143.980 3358.820 144.380 3360.170 ;
        RECT 144.680 3356.270 145.080 3360.170 ;
        RECT 142.230 3355.470 142.680 3355.920 ;
        RECT 145.330 3355.470 145.780 3355.920 ;
        RECT 143.180 3352.270 143.580 3355.170 ;
        RECT 143.980 3352.270 144.380 3353.620 ;
        RECT 144.680 3352.270 145.080 3355.170 ;
        RECT 146.280 3353.170 146.680 3359.270 ;
        RECT 147.880 3356.270 148.280 3360.170 ;
        RECT 148.680 3359.220 149.080 3360.170 ;
        RECT 149.380 3359.220 149.780 3359.270 ;
        RECT 148.680 3358.720 149.780 3359.220 ;
        RECT 149.380 3356.270 149.780 3358.720 ;
        RECT 150.980 3355.970 151.380 3359.270 ;
        RECT 151.780 3359.220 152.180 3360.170 ;
        RECT 152.480 3359.220 152.880 3359.270 ;
        RECT 151.780 3358.720 152.880 3359.220 ;
        RECT 152.480 3356.270 152.880 3358.720 ;
        RECT 146.930 3355.470 147.380 3355.920 ;
        RECT 149.780 3355.470 150.730 3355.970 ;
        RECT 150.980 3355.470 153.830 3355.970 ;
        RECT 147.880 3352.270 148.280 3355.170 ;
        RECT 149.380 3353.620 149.780 3355.170 ;
        RECT 148.680 3353.170 149.780 3353.620 ;
        RECT 150.980 3353.170 151.380 3355.470 ;
        RECT 152.480 3353.620 152.880 3355.170 ;
        RECT 151.780 3353.170 152.880 3353.620 ;
        RECT 154.080 3353.170 154.480 3359.270 ;
        RECT 154.880 3358.820 155.280 3360.170 ;
        RECT 155.580 3356.270 155.980 3360.170 ;
        RECT 156.230 3355.470 156.680 3355.920 ;
        RECT 148.680 3353.120 149.080 3353.170 ;
        RECT 149.380 3352.270 149.780 3353.170 ;
        RECT 151.780 3353.120 152.180 3353.170 ;
        RECT 152.480 3352.270 152.880 3353.170 ;
        RECT 154.880 3352.270 155.280 3353.620 ;
        RECT 155.580 3352.270 155.980 3355.170 ;
        RECT 157.180 3353.170 157.580 3359.270 ;
        RECT 158.780 3356.270 159.180 3360.170 ;
        RECT 157.830 3355.470 158.280 3355.920 ;
        RECT 158.780 3352.270 159.180 3355.170 ;
        RECT 112.780 3351.870 159.180 3352.270 ;
        RECT 70.330 3350.775 77.480 3350.790 ;
        RECT 69.120 3350.605 77.480 3350.775 ;
        RECT 68.430 3349.990 68.830 3350.490 ;
        RECT 69.245 3349.465 69.475 3350.605 ;
        RECT 70.145 3350.440 77.480 3350.605 ;
        RECT 69.645 3349.455 69.975 3350.435 ;
        RECT 70.145 3349.465 70.355 3350.440 ;
        RECT 77.130 3350.305 77.480 3350.440 ;
        RECT 77.130 3350.135 80.350 3350.305 ;
        RECT 81.710 3350.290 83.550 3350.305 ;
        RECT 87.830 3350.290 88.180 3350.740 ;
        RECT 81.710 3350.135 88.180 3350.290 ;
        RECT 69.225 3349.045 69.555 3349.295 ;
        RECT 69.725 3349.240 69.975 3349.455 ;
        RECT 77.215 3349.285 77.595 3349.965 ;
        RECT 78.185 3349.285 78.355 3350.135 ;
        RECT 78.525 3349.455 78.855 3349.965 ;
        RECT 79.025 3349.625 79.195 3350.135 ;
        RECT 79.365 3349.455 79.765 3349.965 ;
        RECT 78.525 3349.285 79.765 3349.455 ;
        RECT 69.725 3349.070 69.980 3349.240 ;
        RECT 68.430 3348.240 68.830 3348.740 ;
        RECT 69.245 3348.055 69.475 3348.875 ;
        RECT 69.725 3348.855 69.975 3349.070 ;
        RECT 69.645 3348.225 69.975 3348.855 ;
        RECT 70.145 3348.240 70.355 3348.875 ;
        RECT 77.215 3348.325 77.385 3349.285 ;
        RECT 77.555 3348.945 78.860 3349.115 ;
        RECT 79.945 3349.035 80.265 3349.965 ;
        RECT 80.880 3349.240 81.280 3349.740 ;
        RECT 81.885 3349.205 82.055 3349.965 ;
        RECT 82.270 3349.375 82.600 3350.135 ;
        RECT 81.885 3349.035 82.600 3349.205 ;
        RECT 82.770 3349.060 83.025 3349.965 ;
        RECT 77.555 3348.495 77.800 3348.945 ;
        RECT 77.970 3348.575 78.520 3348.775 ;
        RECT 78.690 3348.745 78.860 3348.945 ;
        RECT 79.635 3348.890 80.265 3349.035 ;
        RECT 79.635 3348.840 81.480 3348.890 ;
        RECT 81.795 3348.840 82.150 3348.855 ;
        RECT 78.690 3348.575 79.065 3348.745 ;
        RECT 79.235 3348.325 79.465 3348.825 ;
        RECT 70.145 3348.055 75.030 3348.240 ;
        RECT 77.215 3348.155 79.465 3348.325 ;
        RECT 79.635 3348.640 82.150 3348.840 ;
        RECT 69.120 3347.890 75.030 3348.055 ;
        RECT 69.120 3347.885 70.500 3347.890 ;
        RECT 74.680 3347.690 75.030 3347.890 ;
        RECT 77.265 3347.690 77.595 3347.975 ;
        RECT 77.765 3347.835 77.935 3348.155 ;
        RECT 79.635 3347.985 79.805 3348.640 ;
        RECT 81.795 3348.485 82.150 3348.640 ;
        RECT 82.430 3348.825 82.600 3349.035 ;
        RECT 82.430 3348.495 82.685 3348.825 ;
        RECT 74.680 3347.585 77.595 3347.690 ;
        RECT 78.105 3347.585 78.435 3347.975 ;
        RECT 78.850 3347.815 79.805 3347.985 ;
        RECT 79.975 3347.585 80.265 3348.420 ;
        RECT 82.430 3348.305 82.600 3348.495 ;
        RECT 82.855 3348.330 83.025 3349.060 ;
        RECT 83.200 3349.940 88.180 3350.135 ;
        RECT 108.080 3350.470 108.680 3350.920 ;
        RECT 108.080 3349.970 114.080 3350.470 ;
        RECT 83.200 3348.985 83.460 3349.940 ;
        RECT 87.830 3349.540 88.180 3349.940 ;
        RECT 83.830 3348.520 108.730 3348.920 ;
        RECT 80.780 3347.740 81.280 3348.140 ;
        RECT 81.885 3348.135 82.600 3348.305 ;
        RECT 81.885 3347.755 82.055 3348.135 ;
        RECT 82.270 3347.585 82.600 3347.965 ;
        RECT 82.770 3347.755 83.025 3348.330 ;
        RECT 83.200 3347.585 83.460 3348.425 ;
        RECT 108.330 3348.120 108.730 3348.520 ;
        RECT 113.580 3348.370 114.080 3349.970 ;
        RECT 120.620 3349.495 122.920 3349.665 ;
        RECT 119.980 3348.650 120.280 3349.150 ;
        RECT 120.705 3348.925 120.965 3349.325 ;
        RECT 121.135 3349.095 122.070 3349.495 ;
        RECT 122.240 3349.320 122.835 3349.325 ;
        RECT 122.240 3349.020 125.130 3349.320 ;
        RECT 122.240 3348.985 122.835 3349.020 ;
        RECT 120.705 3348.755 122.070 3348.925 ;
        RECT 113.580 3347.820 114.780 3348.370 ;
        RECT 120.705 3347.855 121.165 3348.585 ;
        RECT 121.335 3347.685 122.070 3348.755 ;
        RECT 74.680 3347.415 80.350 3347.585 ;
        RECT 81.710 3347.415 83.550 3347.585 ;
        RECT 74.680 3347.340 77.330 3347.415 ;
        RECT 71.230 3345.615 72.530 3345.740 ;
        RECT 74.680 3345.615 75.030 3347.340 ;
        RECT 120.030 3347.020 120.380 3347.570 ;
        RECT 120.705 3347.515 122.070 3347.685 ;
        RECT 122.240 3347.665 122.415 3348.985 ;
        RECT 122.595 3348.170 122.835 3348.815 ;
        RECT 122.595 3347.870 122.980 3348.170 ;
        RECT 122.595 3347.835 122.835 3347.870 ;
        RECT 120.705 3347.115 120.965 3347.515 ;
        RECT 121.135 3346.945 122.070 3347.345 ;
        RECT 122.240 3347.115 122.835 3347.665 ;
        RECT 120.620 3346.775 122.920 3346.945 ;
        RECT 124.830 3346.170 125.130 3349.020 ;
        RECT 127.230 3348.270 127.630 3351.870 ;
        RECT 157.630 3348.370 158.030 3351.870 ;
        RECT 157.630 3348.270 171.230 3348.370 ;
        RECT 127.230 3347.870 171.230 3348.270 ;
        RECT 82.080 3345.615 84.230 3345.640 ;
        RECT 85.530 3345.615 91.880 3345.970 ;
        RECT 124.780 3345.770 125.180 3346.170 ;
        RECT 69.980 3345.470 91.880 3345.615 ;
        RECT 69.980 3345.445 85.880 3345.470 ;
        RECT 70.125 3344.625 70.335 3345.445 ;
        RECT 71.005 3345.290 72.530 3345.445 ;
        RECT 70.505 3344.645 70.835 3345.275 ;
        RECT 70.505 3344.045 70.755 3344.645 ;
        RECT 71.005 3344.625 71.235 3345.290 ;
        RECT 72.910 3344.735 73.165 3345.265 ;
        RECT 73.345 3344.985 73.630 3345.445 ;
        RECT 70.925 3344.450 71.255 3344.455 ;
        RECT 72.910 3344.450 73.090 3344.735 ;
        RECT 73.810 3344.535 74.060 3345.185 ;
        RECT 70.925 3344.210 73.090 3344.450 ;
        RECT 70.925 3344.205 71.255 3344.210 ;
        RECT 70.125 3342.895 70.335 3344.035 ;
        RECT 70.505 3343.065 70.835 3344.045 ;
        RECT 71.005 3342.895 71.235 3344.035 ;
        RECT 72.910 3343.875 73.090 3344.210 ;
        RECT 73.260 3344.205 74.060 3344.535 ;
        RECT 71.830 3343.290 72.230 3343.790 ;
        RECT 72.910 3343.205 73.165 3343.875 ;
        RECT 73.345 3342.895 73.630 3343.695 ;
        RECT 73.810 3343.615 74.060 3344.205 ;
        RECT 74.260 3344.850 74.580 3345.180 ;
        RECT 74.760 3344.965 75.420 3345.445 ;
        RECT 75.620 3345.055 76.470 3345.225 ;
        RECT 74.260 3343.955 74.450 3344.850 ;
        RECT 74.770 3344.525 75.430 3344.795 ;
        RECT 75.100 3344.465 75.430 3344.525 ;
        RECT 74.620 3344.295 74.950 3344.355 ;
        RECT 75.620 3344.295 75.790 3345.055 ;
        RECT 77.030 3344.985 77.350 3345.445 ;
        RECT 77.550 3344.805 77.800 3345.235 ;
        RECT 78.090 3345.005 78.500 3345.445 ;
        RECT 78.670 3345.065 79.685 3345.265 ;
        RECT 75.960 3344.635 77.210 3344.805 ;
        RECT 75.960 3344.515 76.290 3344.635 ;
        RECT 74.620 3344.125 76.520 3344.295 ;
        RECT 74.260 3343.785 76.180 3343.955 ;
        RECT 74.260 3343.765 74.580 3343.785 ;
        RECT 73.810 3343.105 74.140 3343.615 ;
        RECT 74.410 3343.155 74.580 3343.765 ;
        RECT 76.350 3343.615 76.520 3344.125 ;
        RECT 76.690 3344.055 76.870 3344.465 ;
        RECT 77.040 3343.875 77.210 3344.635 ;
        RECT 74.750 3342.895 75.080 3343.585 ;
        RECT 75.310 3343.445 76.520 3343.615 ;
        RECT 76.690 3343.565 77.210 3343.875 ;
        RECT 77.380 3344.465 77.800 3344.805 ;
        RECT 78.090 3344.465 78.500 3344.795 ;
        RECT 77.380 3343.695 77.570 3344.465 ;
        RECT 78.670 3344.335 78.840 3345.065 ;
        RECT 79.985 3344.895 80.155 3345.225 ;
        RECT 80.325 3345.065 80.655 3345.445 ;
        RECT 79.010 3344.515 79.360 3344.885 ;
        RECT 78.670 3344.295 79.090 3344.335 ;
        RECT 77.740 3344.125 79.090 3344.295 ;
        RECT 77.740 3343.965 77.990 3344.125 ;
        RECT 78.500 3343.695 78.750 3343.955 ;
        RECT 77.380 3343.445 78.750 3343.695 ;
        RECT 75.310 3343.155 75.550 3343.445 ;
        RECT 76.350 3343.365 76.520 3343.445 ;
        RECT 75.750 3342.895 76.170 3343.275 ;
        RECT 76.350 3343.115 76.980 3343.365 ;
        RECT 77.450 3342.895 77.780 3343.275 ;
        RECT 77.950 3343.155 78.120 3343.445 ;
        RECT 78.920 3343.280 79.090 3344.125 ;
        RECT 79.540 3343.955 79.760 3344.825 ;
        RECT 79.985 3344.705 80.680 3344.895 ;
        RECT 79.260 3343.575 79.760 3343.955 ;
        RECT 79.930 3343.905 80.340 3344.525 ;
        RECT 80.510 3343.735 80.680 3344.705 ;
        RECT 79.985 3343.565 80.680 3343.735 ;
        RECT 78.300 3342.895 78.680 3343.275 ;
        RECT 78.920 3343.110 79.750 3343.280 ;
        RECT 79.985 3343.065 80.155 3343.565 ;
        RECT 80.325 3342.895 80.655 3343.395 ;
        RECT 80.870 3343.065 81.095 3345.185 ;
        RECT 81.265 3345.065 81.595 3345.445 ;
        RECT 82.080 3345.290 84.390 3345.445 ;
        RECT 81.765 3344.895 81.935 3345.185 ;
        RECT 81.270 3344.725 81.935 3344.895 ;
        RECT 83.180 3344.890 83.680 3345.290 ;
        RECT 81.270 3343.735 81.500 3344.725 ;
        RECT 84.130 3344.605 84.390 3345.290 ;
        RECT 84.565 3344.700 84.820 3345.275 ;
        RECT 84.990 3345.065 85.320 3345.445 ;
        RECT 85.535 3344.895 85.705 3345.275 ;
        RECT 127.230 3344.970 127.630 3347.870 ;
        RECT 84.990 3344.725 85.705 3344.895 ;
        RECT 81.670 3344.540 82.020 3344.555 ;
        RECT 81.670 3344.190 83.580 3344.540 ;
        RECT 81.670 3343.905 82.020 3344.190 ;
        RECT 81.270 3343.565 81.935 3343.735 ;
        RECT 81.265 3342.895 81.595 3343.395 ;
        RECT 81.765 3343.065 81.935 3343.565 ;
        RECT 84.130 3342.895 84.390 3344.045 ;
        RECT 84.565 3343.970 84.735 3344.700 ;
        RECT 84.990 3344.535 85.160 3344.725 ;
        RECT 86.080 3344.550 98.780 3344.720 ;
        RECT 84.905 3344.205 85.160 3344.535 ;
        RECT 84.990 3343.995 85.160 3344.205 ;
        RECT 85.440 3344.170 98.780 3344.550 ;
        RECT 128.130 3344.220 128.580 3344.670 ;
        RECT 86.080 3344.120 98.780 3344.170 ;
        RECT 84.565 3343.065 84.820 3343.970 ;
        RECT 84.990 3343.825 85.705 3343.995 ;
        RECT 84.990 3342.895 85.320 3343.655 ;
        RECT 85.535 3343.065 85.705 3343.825 ;
        RECT 98.180 3343.520 98.780 3344.120 ;
        RECT 87.830 3342.940 88.180 3343.390 ;
        RECT 85.830 3342.895 88.180 3342.940 ;
        RECT 69.980 3342.725 71.360 3342.895 ;
        RECT 72.450 3342.725 82.110 3342.895 ;
        RECT 84.040 3342.725 88.180 3342.895 ;
        RECT 85.830 3342.590 88.180 3342.725 ;
        RECT 127.230 3339.970 127.630 3343.870 ;
        RECT 128.830 3340.870 129.230 3346.970 ;
        RECT 130.430 3344.970 130.830 3347.870 ;
        RECT 131.130 3346.520 131.530 3347.870 ;
        RECT 133.530 3346.970 133.930 3347.870 ;
        RECT 134.230 3346.970 134.630 3347.020 ;
        RECT 136.630 3346.970 137.030 3347.870 ;
        RECT 137.330 3346.970 137.730 3347.020 ;
        RECT 129.730 3344.220 130.180 3344.670 ;
        RECT 130.430 3339.970 130.830 3343.870 ;
        RECT 131.130 3339.970 131.530 3341.320 ;
        RECT 131.930 3340.870 132.330 3346.970 ;
        RECT 133.530 3346.520 134.630 3346.970 ;
        RECT 133.530 3344.970 133.930 3346.520 ;
        RECT 135.030 3344.670 135.430 3346.970 ;
        RECT 136.630 3346.520 137.730 3346.970 ;
        RECT 136.630 3344.970 137.030 3346.520 ;
        RECT 138.130 3344.970 138.530 3347.870 ;
        RECT 132.580 3344.170 135.430 3344.670 ;
        RECT 135.680 3344.170 136.630 3344.670 ;
        RECT 139.030 3344.220 139.480 3344.670 ;
        RECT 133.530 3341.420 133.930 3343.870 ;
        RECT 133.530 3340.920 134.630 3341.420 ;
        RECT 133.530 3340.870 133.930 3340.920 ;
        RECT 134.230 3339.970 134.630 3340.920 ;
        RECT 135.030 3340.870 135.430 3344.170 ;
        RECT 136.630 3341.420 137.030 3343.870 ;
        RECT 136.630 3340.920 137.730 3341.420 ;
        RECT 136.630 3340.870 137.030 3340.920 ;
        RECT 137.330 3339.970 137.730 3340.920 ;
        RECT 138.130 3339.970 138.530 3343.870 ;
        RECT 139.730 3340.870 140.130 3346.970 ;
        RECT 141.330 3344.970 141.730 3347.870 ;
        RECT 142.030 3346.520 142.430 3347.870 ;
        RECT 142.830 3344.970 143.230 3347.870 ;
        RECT 140.630 3344.220 141.080 3344.670 ;
        RECT 143.730 3344.220 144.180 3344.670 ;
        RECT 141.330 3339.970 141.730 3343.870 ;
        RECT 142.030 3339.970 142.430 3341.320 ;
        RECT 142.830 3339.970 143.230 3343.870 ;
        RECT 144.430 3340.870 144.830 3346.970 ;
        RECT 146.030 3344.970 146.430 3347.870 ;
        RECT 146.730 3346.520 147.130 3347.870 ;
        RECT 149.130 3346.970 149.530 3347.870 ;
        RECT 149.830 3346.970 150.230 3347.020 ;
        RECT 152.230 3346.970 152.630 3347.870 ;
        RECT 152.930 3346.970 153.330 3347.020 ;
        RECT 145.330 3344.220 145.780 3344.670 ;
        RECT 146.030 3339.970 146.430 3343.870 ;
        RECT 146.730 3339.970 147.130 3341.320 ;
        RECT 147.530 3340.870 147.930 3346.970 ;
        RECT 149.130 3346.520 150.230 3346.970 ;
        RECT 149.130 3344.970 149.530 3346.520 ;
        RECT 150.630 3344.670 151.030 3346.970 ;
        RECT 152.230 3346.520 153.330 3346.970 ;
        RECT 152.230 3344.970 152.630 3346.520 ;
        RECT 153.730 3344.970 154.130 3347.870 ;
        RECT 148.180 3344.170 151.030 3344.670 ;
        RECT 151.280 3344.170 152.230 3344.670 ;
        RECT 154.630 3344.220 155.080 3344.670 ;
        RECT 149.130 3341.420 149.530 3343.870 ;
        RECT 149.130 3340.920 150.230 3341.420 ;
        RECT 149.130 3340.870 149.530 3340.920 ;
        RECT 149.830 3339.970 150.230 3340.920 ;
        RECT 150.630 3340.870 151.030 3344.170 ;
        RECT 152.230 3341.420 152.630 3343.870 ;
        RECT 152.230 3340.920 153.330 3341.420 ;
        RECT 152.230 3340.870 152.630 3340.920 ;
        RECT 152.930 3339.970 153.330 3340.920 ;
        RECT 153.730 3339.970 154.130 3343.870 ;
        RECT 155.330 3340.870 155.730 3346.970 ;
        RECT 156.930 3344.970 157.330 3347.870 ;
        RECT 157.630 3346.520 158.030 3347.870 ;
        RECT 170.730 3347.270 171.230 3347.870 ;
        RECT 156.230 3344.220 156.680 3344.670 ;
        RECT 156.930 3339.970 157.330 3343.870 ;
        RECT 157.630 3339.970 158.030 3341.320 ;
        RECT 127.230 3339.570 158.030 3339.970 ;
        RECT 70.780 3336.965 71.180 3337.120 ;
        RECT 70.770 3336.795 74.450 3336.965 ;
        RECT 74.870 3336.795 78.550 3336.965 ;
        RECT 78.970 3336.795 82.650 3336.965 ;
        RECT 83.370 3336.795 87.050 3336.965 ;
        RECT 87.470 3336.795 91.150 3336.965 ;
        RECT 91.570 3336.795 95.250 3336.965 ;
        RECT 70.970 3336.165 71.255 3336.625 ;
        RECT 71.425 3336.335 71.695 3336.795 ;
        RECT 70.970 3335.945 71.925 3336.165 ;
        RECT 70.855 3335.215 71.545 3335.775 ;
        RECT 71.715 3335.045 71.925 3335.945 ;
        RECT 70.970 3334.875 71.925 3335.045 ;
        RECT 72.095 3335.775 72.495 3336.625 ;
        RECT 72.685 3336.165 72.965 3336.625 ;
        RECT 73.485 3336.335 73.810 3336.795 ;
        RECT 72.685 3335.945 73.810 3336.165 ;
        RECT 72.095 3335.215 73.190 3335.775 ;
        RECT 73.360 3335.485 73.810 3335.945 ;
        RECT 73.980 3335.770 74.365 3336.625 ;
        RECT 75.070 3336.165 75.355 3336.625 ;
        RECT 75.525 3336.335 75.795 3336.795 ;
        RECT 75.070 3335.945 76.025 3336.165 ;
        RECT 74.955 3335.770 75.645 3335.775 ;
        RECT 73.980 3335.655 75.645 3335.770 ;
        RECT 70.970 3334.415 71.255 3334.875 ;
        RECT 71.425 3334.245 71.695 3334.705 ;
        RECT 72.095 3334.415 72.495 3335.215 ;
        RECT 73.360 3335.155 73.915 3335.485 ;
        RECT 74.085 3335.220 75.645 3335.655 ;
        RECT 73.360 3335.045 73.810 3335.155 ;
        RECT 72.685 3334.875 73.810 3335.045 ;
        RECT 74.085 3334.985 74.365 3335.220 ;
        RECT 74.955 3335.215 75.645 3335.220 ;
        RECT 75.815 3335.045 76.025 3335.945 ;
        RECT 72.685 3334.415 72.965 3334.875 ;
        RECT 73.485 3334.245 73.810 3334.705 ;
        RECT 73.980 3334.415 74.365 3334.985 ;
        RECT 75.070 3334.875 76.025 3335.045 ;
        RECT 76.195 3335.775 76.595 3336.625 ;
        RECT 76.785 3336.165 77.065 3336.625 ;
        RECT 77.585 3336.335 77.910 3336.795 ;
        RECT 76.785 3335.945 77.910 3336.165 ;
        RECT 76.195 3335.215 77.290 3335.775 ;
        RECT 77.460 3335.485 77.910 3335.945 ;
        RECT 78.080 3335.770 78.465 3336.625 ;
        RECT 79.170 3336.165 79.455 3336.625 ;
        RECT 79.625 3336.335 79.895 3336.795 ;
        RECT 79.170 3335.945 80.125 3336.165 ;
        RECT 79.055 3335.770 79.745 3335.775 ;
        RECT 78.080 3335.655 79.745 3335.770 ;
        RECT 75.070 3334.415 75.355 3334.875 ;
        RECT 75.525 3334.245 75.795 3334.705 ;
        RECT 76.195 3334.415 76.595 3335.215 ;
        RECT 77.460 3335.155 78.015 3335.485 ;
        RECT 78.185 3335.220 79.745 3335.655 ;
        RECT 77.460 3335.045 77.910 3335.155 ;
        RECT 76.785 3334.875 77.910 3335.045 ;
        RECT 78.185 3334.985 78.465 3335.220 ;
        RECT 79.055 3335.215 79.745 3335.220 ;
        RECT 79.915 3335.045 80.125 3335.945 ;
        RECT 76.785 3334.415 77.065 3334.875 ;
        RECT 77.585 3334.245 77.910 3334.705 ;
        RECT 78.080 3334.415 78.465 3334.985 ;
        RECT 79.170 3334.875 80.125 3335.045 ;
        RECT 80.295 3335.775 80.695 3336.625 ;
        RECT 80.885 3336.165 81.165 3336.625 ;
        RECT 81.685 3336.335 82.010 3336.795 ;
        RECT 80.885 3335.945 82.010 3336.165 ;
        RECT 80.295 3335.215 81.390 3335.775 ;
        RECT 81.560 3335.485 82.010 3335.945 ;
        RECT 82.180 3335.770 82.565 3336.625 ;
        RECT 82.880 3335.970 83.280 3336.470 ;
        RECT 83.570 3336.165 83.855 3336.625 ;
        RECT 84.025 3336.335 84.295 3336.795 ;
        RECT 83.570 3335.945 84.525 3336.165 ;
        RECT 83.455 3335.770 84.145 3335.775 ;
        RECT 82.180 3335.655 84.145 3335.770 ;
        RECT 79.170 3334.415 79.455 3334.875 ;
        RECT 79.625 3334.245 79.895 3334.705 ;
        RECT 80.295 3334.415 80.695 3335.215 ;
        RECT 81.560 3335.155 82.115 3335.485 ;
        RECT 82.285 3335.220 84.145 3335.655 ;
        RECT 81.560 3335.045 82.010 3335.155 ;
        RECT 80.885 3334.875 82.010 3335.045 ;
        RECT 82.285 3334.985 82.565 3335.220 ;
        RECT 83.455 3335.215 84.145 3335.220 ;
        RECT 84.315 3335.045 84.525 3335.945 ;
        RECT 80.885 3334.415 81.165 3334.875 ;
        RECT 81.685 3334.245 82.010 3334.705 ;
        RECT 82.180 3334.415 82.565 3334.985 ;
        RECT 82.830 3334.410 83.140 3334.910 ;
        RECT 83.570 3334.875 84.525 3335.045 ;
        RECT 84.695 3335.775 85.095 3336.625 ;
        RECT 85.285 3336.165 85.565 3336.625 ;
        RECT 86.085 3336.335 86.410 3336.795 ;
        RECT 85.285 3335.945 86.410 3336.165 ;
        RECT 84.695 3335.215 85.790 3335.775 ;
        RECT 85.960 3335.485 86.410 3335.945 ;
        RECT 86.580 3335.770 86.965 3336.625 ;
        RECT 87.670 3336.165 87.955 3336.625 ;
        RECT 88.125 3336.335 88.395 3336.795 ;
        RECT 87.670 3335.945 88.625 3336.165 ;
        RECT 87.555 3335.770 88.245 3335.775 ;
        RECT 86.580 3335.655 88.245 3335.770 ;
        RECT 83.570 3334.415 83.855 3334.875 ;
        RECT 84.025 3334.245 84.295 3334.705 ;
        RECT 84.695 3334.415 85.095 3335.215 ;
        RECT 85.960 3335.155 86.515 3335.485 ;
        RECT 86.685 3335.220 88.245 3335.655 ;
        RECT 85.960 3335.045 86.410 3335.155 ;
        RECT 85.285 3334.875 86.410 3335.045 ;
        RECT 86.685 3334.985 86.965 3335.220 ;
        RECT 87.555 3335.215 88.245 3335.220 ;
        RECT 88.415 3335.045 88.625 3335.945 ;
        RECT 85.285 3334.415 85.565 3334.875 ;
        RECT 86.085 3334.245 86.410 3334.705 ;
        RECT 86.580 3334.415 86.965 3334.985 ;
        RECT 87.670 3334.875 88.625 3335.045 ;
        RECT 88.795 3335.775 89.195 3336.625 ;
        RECT 89.385 3336.165 89.665 3336.625 ;
        RECT 90.185 3336.335 90.510 3336.795 ;
        RECT 89.385 3335.945 90.510 3336.165 ;
        RECT 88.795 3335.215 89.890 3335.775 ;
        RECT 90.060 3335.485 90.510 3335.945 ;
        RECT 90.680 3335.770 91.065 3336.625 ;
        RECT 91.770 3336.165 92.055 3336.625 ;
        RECT 92.225 3336.335 92.495 3336.795 ;
        RECT 91.770 3335.945 92.725 3336.165 ;
        RECT 91.655 3335.770 92.345 3335.775 ;
        RECT 90.680 3335.655 92.345 3335.770 ;
        RECT 87.670 3334.415 87.955 3334.875 ;
        RECT 88.125 3334.245 88.395 3334.705 ;
        RECT 88.795 3334.415 89.195 3335.215 ;
        RECT 90.060 3335.155 90.615 3335.485 ;
        RECT 90.785 3335.220 92.345 3335.655 ;
        RECT 90.060 3335.045 90.510 3335.155 ;
        RECT 89.385 3334.875 90.510 3335.045 ;
        RECT 90.785 3334.985 91.065 3335.220 ;
        RECT 91.655 3335.215 92.345 3335.220 ;
        RECT 92.515 3335.045 92.725 3335.945 ;
        RECT 89.385 3334.415 89.665 3334.875 ;
        RECT 90.185 3334.245 90.510 3334.705 ;
        RECT 90.680 3334.415 91.065 3334.985 ;
        RECT 91.770 3334.875 92.725 3335.045 ;
        RECT 92.895 3335.775 93.295 3336.625 ;
        RECT 93.485 3336.165 93.765 3336.625 ;
        RECT 94.285 3336.335 94.610 3336.795 ;
        RECT 93.485 3335.945 94.610 3336.165 ;
        RECT 92.895 3335.215 93.990 3335.775 ;
        RECT 94.160 3335.485 94.610 3335.945 ;
        RECT 94.780 3335.655 95.165 3336.625 ;
        RECT 91.770 3334.415 92.055 3334.875 ;
        RECT 92.225 3334.245 92.495 3334.705 ;
        RECT 92.895 3334.415 93.295 3335.215 ;
        RECT 94.160 3335.155 94.715 3335.485 ;
        RECT 94.160 3335.045 94.610 3335.155 ;
        RECT 93.485 3334.875 94.610 3335.045 ;
        RECT 94.885 3335.070 95.165 3335.655 ;
        RECT 94.885 3334.985 96.580 3335.070 ;
        RECT 93.485 3334.415 93.765 3334.875 ;
        RECT 94.780 3334.720 96.580 3334.985 ;
        RECT 94.285 3334.245 94.610 3334.705 ;
        RECT 94.780 3334.415 95.165 3334.720 ;
        RECT 70.770 3334.075 74.450 3334.245 ;
        RECT 74.870 3334.075 78.550 3334.245 ;
        RECT 78.970 3334.075 82.650 3334.245 ;
        RECT 83.370 3334.075 87.050 3334.245 ;
        RECT 87.470 3334.075 91.150 3334.245 ;
        RECT 91.570 3334.075 95.250 3334.245 ;
        RECT 96.230 3333.720 96.580 3334.720 ;
        RECT 85.630 3333.370 96.580 3333.720 ;
        RECT 72.230 3332.965 74.980 3333.120 ;
        RECT 70.770 3332.920 81.930 3332.965 ;
        RECT 70.770 3332.795 72.610 3332.920 ;
        RECT 70.945 3331.865 71.115 3332.625 ;
        RECT 71.330 3332.035 71.660 3332.795 ;
        RECT 70.945 3331.695 71.660 3331.865 ;
        RECT 71.830 3331.720 72.085 3332.625 ;
        RECT 70.855 3331.145 71.210 3331.515 ;
        RECT 71.490 3331.485 71.660 3331.695 ;
        RECT 71.490 3331.155 71.745 3331.485 ;
        RECT 71.490 3330.965 71.660 3331.155 ;
        RECT 71.915 3330.990 72.085 3331.720 ;
        RECT 72.260 3331.645 72.520 3332.795 ;
        RECT 73.030 3331.970 73.430 3332.920 ;
        RECT 74.570 3332.795 81.930 3332.920 ;
        RECT 83.820 3332.795 85.200 3332.965 ;
        RECT 74.745 3332.125 74.915 3332.625 ;
        RECT 75.085 3332.295 75.415 3332.795 ;
        RECT 74.745 3331.955 75.410 3332.125 ;
        RECT 74.660 3331.135 75.010 3331.785 ;
        RECT 70.945 3330.795 71.660 3330.965 ;
        RECT 70.945 3330.415 71.115 3330.795 ;
        RECT 71.330 3330.245 71.660 3330.625 ;
        RECT 71.830 3330.415 72.085 3330.990 ;
        RECT 72.260 3330.245 72.520 3331.085 ;
        RECT 72.780 3330.520 73.180 3331.020 ;
        RECT 75.180 3330.965 75.410 3331.955 ;
        RECT 74.745 3330.795 75.410 3330.965 ;
        RECT 74.745 3330.505 74.915 3330.795 ;
        RECT 75.085 3330.245 75.415 3330.625 ;
        RECT 75.585 3330.505 75.770 3332.625 ;
        RECT 76.010 3332.335 76.275 3332.795 ;
        RECT 76.445 3332.200 76.695 3332.625 ;
        RECT 76.905 3332.350 78.010 3332.520 ;
        RECT 76.390 3332.070 76.695 3332.200 ;
        RECT 75.940 3330.875 76.220 3331.825 ;
        RECT 76.390 3330.965 76.560 3332.070 ;
        RECT 76.730 3331.285 76.970 3331.880 ;
        RECT 77.140 3331.815 77.670 3332.180 ;
        RECT 77.140 3331.115 77.310 3331.815 ;
        RECT 77.840 3331.735 78.010 3332.350 ;
        RECT 78.180 3331.995 78.350 3332.795 ;
        RECT 78.520 3332.295 78.770 3332.625 ;
        RECT 78.995 3332.325 79.880 3332.495 ;
        RECT 77.840 3331.645 78.350 3331.735 ;
        RECT 76.390 3330.835 76.615 3330.965 ;
        RECT 76.785 3330.895 77.310 3331.115 ;
        RECT 77.480 3331.475 78.350 3331.645 ;
        RECT 76.025 3330.245 76.275 3330.705 ;
        RECT 76.445 3330.695 76.615 3330.835 ;
        RECT 77.480 3330.695 77.650 3331.475 ;
        RECT 78.180 3331.405 78.350 3331.475 ;
        RECT 77.860 3331.225 78.060 3331.255 ;
        RECT 78.520 3331.225 78.690 3332.295 ;
        RECT 78.860 3331.405 79.050 3332.125 ;
        RECT 77.860 3330.925 78.690 3331.225 ;
        RECT 79.220 3331.195 79.540 3332.155 ;
        RECT 76.445 3330.525 76.780 3330.695 ;
        RECT 76.975 3330.525 77.650 3330.695 ;
        RECT 77.970 3330.245 78.340 3330.745 ;
        RECT 78.520 3330.695 78.690 3330.925 ;
        RECT 79.075 3330.865 79.540 3331.195 ;
        RECT 79.710 3331.485 79.880 3332.325 ;
        RECT 80.060 3332.295 80.375 3332.795 ;
        RECT 80.605 3332.065 80.945 3332.625 ;
        RECT 80.050 3331.690 80.945 3332.065 ;
        RECT 81.115 3331.785 81.285 3332.795 ;
        RECT 80.755 3331.485 80.945 3331.690 ;
        RECT 81.455 3331.735 81.785 3332.580 ;
        RECT 81.455 3331.655 81.845 3331.735 ;
        RECT 83.905 3331.655 84.185 3332.795 ;
        RECT 81.630 3331.605 81.845 3331.655 ;
        RECT 84.355 3331.645 84.685 3332.625 ;
        RECT 84.855 3331.655 85.115 3332.795 ;
        RECT 79.710 3331.155 80.585 3331.485 ;
        RECT 80.755 3331.155 81.505 3331.485 ;
        RECT 81.675 3331.470 81.845 3331.605 ;
        RECT 83.915 3331.470 84.250 3331.485 ;
        RECT 81.675 3331.220 84.250 3331.470 ;
        RECT 79.710 3330.695 79.880 3331.155 ;
        RECT 80.755 3330.985 80.955 3331.155 ;
        RECT 81.675 3331.025 81.845 3331.220 ;
        RECT 81.620 3330.985 81.845 3331.025 ;
        RECT 78.520 3330.525 78.925 3330.695 ;
        RECT 79.095 3330.525 79.880 3330.695 ;
        RECT 80.155 3330.245 80.365 3330.775 ;
        RECT 80.625 3330.460 80.955 3330.985 ;
        RECT 81.465 3330.900 81.845 3330.985 ;
        RECT 81.125 3330.245 81.295 3330.855 ;
        RECT 81.465 3330.465 81.795 3330.900 ;
        RECT 70.770 3330.075 72.610 3330.245 ;
        RECT 74.570 3330.075 81.930 3330.245 ;
        RECT 82.430 3326.070 83.430 3331.220 ;
        RECT 83.915 3331.215 84.250 3331.220 ;
        RECT 84.420 3331.045 84.590 3331.645 ;
        RECT 84.760 3331.470 85.095 3331.485 ;
        RECT 85.630 3331.470 85.980 3333.370 ;
        RECT 86.470 3332.795 87.850 3332.965 ;
        RECT 86.595 3331.655 86.825 3332.795 ;
        RECT 86.995 3331.645 87.325 3332.625 ;
        RECT 87.495 3331.655 87.705 3332.795 ;
        RECT 98.180 3332.320 98.780 3332.920 ;
        RECT 88.480 3331.720 98.780 3332.320 ;
        RECT 84.760 3331.235 85.980 3331.470 ;
        RECT 86.575 3331.235 86.905 3331.485 ;
        RECT 85.080 3331.220 85.980 3331.235 ;
        RECT 83.905 3330.245 84.215 3331.045 ;
        RECT 84.420 3330.415 85.115 3331.045 ;
        RECT 86.595 3330.245 86.825 3331.065 ;
        RECT 87.075 3331.045 87.325 3331.645 ;
        RECT 98.180 3331.120 98.780 3331.720 ;
        RECT 115.780 3332.070 122.430 3332.470 ;
        RECT 86.995 3330.415 87.325 3331.045 ;
        RECT 87.495 3330.245 87.705 3331.065 ;
        RECT 83.820 3330.075 85.200 3330.245 ;
        RECT 86.470 3330.075 87.850 3330.245 ;
        RECT 115.780 3330.070 116.180 3332.070 ;
        RECT 116.480 3328.770 116.880 3332.070 ;
        RECT 117.380 3328.770 117.780 3330.570 ;
        RECT 119.530 3330.120 119.930 3332.070 ;
        RECT 120.230 3328.770 120.630 3330.570 ;
        RECT 121.130 3328.770 121.530 3330.570 ;
        RECT 122.030 3328.770 122.430 3332.070 ;
        RECT 122.930 3328.020 123.330 3330.570 ;
        RECT 125.030 3328.020 125.430 3330.620 ;
        RECT 125.730 3328.020 126.130 3330.570 ;
        RECT 122.930 3327.620 126.130 3328.020 ;
        RECT 126.630 3326.070 127.030 3330.570 ;
        RECT 127.530 3328.770 127.930 3330.570 ;
        RECT 128.430 3328.770 128.830 3330.570 ;
        RECT 130.530 3330.070 130.930 3330.570 ;
        RECT 131.230 3328.720 131.630 3330.520 ;
        RECT 132.130 3329.220 132.530 3330.520 ;
        RECT 134.080 3329.220 134.580 3339.570 ;
        RECT 138.220 3336.220 140.060 3336.265 ;
        RECT 143.980 3336.220 144.430 3337.620 ;
        RECT 138.220 3336.095 144.430 3336.220 ;
        RECT 138.395 3335.165 138.565 3335.925 ;
        RECT 138.780 3335.335 139.110 3336.095 ;
        RECT 138.395 3334.995 139.110 3335.165 ;
        RECT 139.280 3335.020 139.535 3335.925 ;
        RECT 138.305 3334.445 138.660 3334.815 ;
        RECT 138.940 3334.785 139.110 3334.995 ;
        RECT 138.940 3334.455 139.195 3334.785 ;
        RECT 138.940 3334.265 139.110 3334.455 ;
        RECT 139.365 3334.290 139.535 3335.020 ;
        RECT 139.710 3335.870 144.430 3336.095 ;
        RECT 139.710 3334.945 139.970 3335.870 ;
        RECT 140.330 3335.020 140.630 3335.870 ;
        RECT 138.395 3334.095 139.110 3334.265 ;
        RECT 138.395 3333.715 138.565 3334.095 ;
        RECT 138.780 3333.545 139.110 3333.925 ;
        RECT 139.280 3333.715 139.535 3334.290 ;
        RECT 139.710 3333.545 139.970 3334.385 ;
        RECT 140.330 3333.770 140.630 3334.270 ;
        RECT 138.220 3333.375 140.060 3333.545 ;
        RECT 144.030 3331.470 144.430 3335.870 ;
        RECT 157.880 3332.365 159.230 3332.520 ;
        RECT 145.970 3332.195 148.270 3332.365 ;
        RECT 150.570 3332.195 159.230 3332.365 ;
        RECT 146.100 3331.055 146.365 3332.195 ;
        RECT 146.535 3331.225 146.865 3332.025 ;
        RECT 147.035 3331.395 147.205 3332.195 ;
        RECT 147.375 3331.245 147.705 3332.025 ;
        RECT 147.875 3331.735 148.085 3332.195 ;
        RECT 150.745 3331.525 150.915 3332.025 ;
        RECT 151.085 3331.695 151.415 3332.195 ;
        RECT 150.745 3331.355 151.410 3331.525 ;
        RECT 147.375 3331.225 148.140 3331.245 ;
        RECT 146.535 3331.170 148.140 3331.225 ;
        RECT 150.660 3331.170 151.010 3331.185 ;
        RECT 146.535 3331.055 151.010 3331.170 ;
        RECT 146.075 3330.635 147.705 3330.885 ;
        RECT 147.875 3330.770 151.010 3331.055 ;
        RECT 147.875 3330.465 148.140 3330.770 ;
        RECT 150.660 3330.535 151.010 3330.770 ;
        RECT 137.830 3329.820 144.430 3330.320 ;
        RECT 146.535 3330.285 148.140 3330.465 ;
        RECT 151.180 3330.365 151.410 3331.355 ;
        RECT 137.830 3329.320 138.330 3329.820 ;
        RECT 146.100 3329.645 146.365 3330.105 ;
        RECT 146.535 3329.815 146.865 3330.285 ;
        RECT 147.035 3329.645 147.205 3330.105 ;
        RECT 147.375 3329.815 147.705 3330.285 ;
        RECT 147.875 3329.645 148.125 3330.110 ;
        RECT 149.180 3329.870 149.730 3330.320 ;
        RECT 150.745 3330.195 151.410 3330.365 ;
        RECT 150.745 3329.905 150.915 3330.195 ;
        RECT 145.970 3329.475 148.270 3329.645 ;
        RECT 132.130 3328.720 134.580 3329.220 ;
        RECT 149.355 3328.995 149.605 3329.870 ;
        RECT 151.085 3329.645 151.415 3330.025 ;
        RECT 151.585 3329.905 151.770 3332.025 ;
        RECT 152.010 3331.735 152.275 3332.195 ;
        RECT 152.445 3331.600 152.695 3332.025 ;
        RECT 152.905 3331.750 154.010 3331.920 ;
        RECT 152.390 3331.470 152.695 3331.600 ;
        RECT 151.940 3330.275 152.220 3331.225 ;
        RECT 152.390 3330.365 152.560 3331.470 ;
        RECT 152.730 3330.685 152.970 3331.280 ;
        RECT 153.140 3331.215 153.670 3331.580 ;
        RECT 153.140 3330.515 153.310 3331.215 ;
        RECT 153.840 3331.135 154.010 3331.750 ;
        RECT 154.180 3331.395 154.350 3332.195 ;
        RECT 154.520 3331.695 154.770 3332.025 ;
        RECT 154.995 3331.725 155.880 3331.895 ;
        RECT 153.840 3331.045 154.350 3331.135 ;
        RECT 152.390 3330.235 152.615 3330.365 ;
        RECT 152.785 3330.295 153.310 3330.515 ;
        RECT 153.480 3330.875 154.350 3331.045 ;
        RECT 152.025 3329.645 152.275 3330.105 ;
        RECT 152.445 3330.095 152.615 3330.235 ;
        RECT 153.480 3330.095 153.650 3330.875 ;
        RECT 154.180 3330.805 154.350 3330.875 ;
        RECT 153.860 3330.625 154.060 3330.655 ;
        RECT 154.520 3330.625 154.690 3331.695 ;
        RECT 154.860 3330.805 155.050 3331.525 ;
        RECT 153.860 3330.325 154.690 3330.625 ;
        RECT 155.220 3330.595 155.540 3331.555 ;
        RECT 152.445 3329.925 152.780 3330.095 ;
        RECT 152.975 3329.925 153.650 3330.095 ;
        RECT 153.970 3329.645 154.340 3330.145 ;
        RECT 154.520 3330.095 154.690 3330.325 ;
        RECT 155.075 3330.265 155.540 3330.595 ;
        RECT 155.710 3330.885 155.880 3331.725 ;
        RECT 156.060 3331.695 156.375 3332.195 ;
        RECT 156.605 3331.465 156.945 3332.025 ;
        RECT 156.050 3331.090 156.945 3331.465 ;
        RECT 157.115 3331.185 157.285 3332.195 ;
        RECT 157.880 3332.170 159.230 3332.195 ;
        RECT 156.755 3330.885 156.945 3331.090 ;
        RECT 157.455 3331.135 157.785 3331.980 ;
        RECT 157.455 3331.055 157.845 3331.135 ;
        RECT 157.630 3331.005 157.845 3331.055 ;
        RECT 155.710 3330.555 156.585 3330.885 ;
        RECT 156.755 3330.555 157.505 3330.885 ;
        RECT 155.710 3330.095 155.880 3330.555 ;
        RECT 156.755 3330.385 156.955 3330.555 ;
        RECT 157.675 3330.425 157.845 3331.005 ;
        RECT 157.620 3330.385 157.845 3330.425 ;
        RECT 154.520 3329.925 154.925 3330.095 ;
        RECT 155.095 3329.925 155.880 3330.095 ;
        RECT 156.155 3329.645 156.365 3330.175 ;
        RECT 156.625 3329.860 156.955 3330.385 ;
        RECT 157.465 3330.300 157.845 3330.385 ;
        RECT 157.125 3329.645 157.295 3330.255 ;
        RECT 157.465 3329.865 157.795 3330.300 ;
        RECT 150.570 3329.475 157.930 3329.645 ;
        RECT 82.430 3325.070 94.580 3326.070 ;
        RECT 118.530 3325.570 130.380 3326.070 ;
        RECT 118.530 3325.070 119.030 3325.570 ;
        RECT 116.130 3324.570 119.030 3325.070 ;
        RECT 85.630 3324.335 88.180 3324.340 ;
        RECT 68.970 3324.165 70.810 3324.335 ;
        RECT 72.410 3324.165 82.070 3324.335 ;
        RECT 83.880 3324.165 88.180 3324.335 ;
        RECT 69.145 3323.235 69.315 3323.995 ;
        RECT 69.530 3323.405 69.860 3324.165 ;
        RECT 69.145 3323.065 69.860 3323.235 ;
        RECT 70.030 3323.090 70.285 3323.995 ;
        RECT 66.980 3322.890 69.030 3322.920 ;
        RECT 66.980 3322.540 69.430 3322.890 ;
        RECT 69.690 3322.855 69.860 3323.065 ;
        RECT 66.980 3322.520 69.410 3322.540 ;
        RECT 66.980 3322.120 67.380 3322.520 ;
        RECT 69.055 3322.515 69.410 3322.520 ;
        RECT 69.690 3322.525 69.945 3322.855 ;
        RECT 70.115 3322.840 70.285 3323.090 ;
        RECT 70.460 3323.015 70.720 3324.165 ;
        RECT 71.430 3323.390 71.830 3323.890 ;
        RECT 72.585 3323.495 72.755 3323.995 ;
        RECT 72.925 3323.665 73.255 3324.165 ;
        RECT 72.585 3323.325 73.250 3323.495 ;
        RECT 72.500 3322.840 72.850 3323.155 ;
        RECT 70.115 3322.640 72.850 3322.840 ;
        RECT 69.690 3322.335 69.860 3322.525 ;
        RECT 70.115 3322.360 70.285 3322.640 ;
        RECT 72.500 3322.505 72.850 3322.640 ;
        RECT 68.380 3321.790 68.780 3322.290 ;
        RECT 69.145 3322.165 69.860 3322.335 ;
        RECT 69.145 3321.785 69.315 3322.165 ;
        RECT 69.530 3321.615 69.860 3321.995 ;
        RECT 70.030 3321.785 70.285 3322.360 ;
        RECT 70.460 3321.790 70.720 3322.455 ;
        RECT 73.020 3322.335 73.250 3323.325 ;
        RECT 72.585 3322.165 73.250 3322.335 ;
        RECT 72.585 3321.875 72.755 3322.165 ;
        RECT 70.460 3321.615 72.430 3321.790 ;
        RECT 72.925 3321.615 73.255 3321.995 ;
        RECT 73.425 3321.875 73.650 3323.995 ;
        RECT 73.865 3323.665 74.195 3324.165 ;
        RECT 74.365 3323.495 74.535 3323.995 ;
        RECT 74.770 3323.780 75.600 3323.950 ;
        RECT 75.840 3323.785 76.220 3324.165 ;
        RECT 73.840 3323.325 74.535 3323.495 ;
        RECT 73.840 3322.355 74.010 3323.325 ;
        RECT 74.180 3322.535 74.590 3323.155 ;
        RECT 74.760 3323.105 75.260 3323.485 ;
        RECT 73.840 3322.165 74.535 3322.355 ;
        RECT 74.760 3322.235 74.980 3323.105 ;
        RECT 75.430 3322.935 75.600 3323.780 ;
        RECT 76.400 3323.615 76.570 3323.905 ;
        RECT 76.740 3323.785 77.070 3324.165 ;
        RECT 77.540 3323.695 78.170 3323.945 ;
        RECT 78.350 3323.785 78.770 3324.165 ;
        RECT 78.000 3323.615 78.170 3323.695 ;
        RECT 78.970 3323.615 79.210 3323.905 ;
        RECT 75.770 3323.365 77.140 3323.615 ;
        RECT 75.770 3323.105 76.020 3323.365 ;
        RECT 76.530 3322.935 76.780 3323.095 ;
        RECT 75.430 3322.765 76.780 3322.935 ;
        RECT 75.430 3322.725 75.850 3322.765 ;
        RECT 75.160 3322.175 75.510 3322.545 ;
        RECT 73.865 3321.615 74.195 3321.995 ;
        RECT 74.365 3321.835 74.535 3322.165 ;
        RECT 75.680 3321.995 75.850 3322.725 ;
        RECT 76.950 3322.595 77.140 3323.365 ;
        RECT 76.020 3322.265 76.430 3322.595 ;
        RECT 76.720 3322.255 77.140 3322.595 ;
        RECT 77.310 3323.185 77.830 3323.495 ;
        RECT 78.000 3323.445 79.210 3323.615 ;
        RECT 79.440 3323.475 79.770 3324.165 ;
        RECT 77.310 3322.425 77.480 3323.185 ;
        RECT 77.650 3322.595 77.830 3323.005 ;
        RECT 78.000 3322.935 78.170 3323.445 ;
        RECT 79.940 3323.295 80.110 3323.905 ;
        RECT 80.380 3323.445 80.710 3323.955 ;
        RECT 79.940 3323.275 80.260 3323.295 ;
        RECT 78.340 3323.105 80.260 3323.275 ;
        RECT 78.000 3322.765 79.900 3322.935 ;
        RECT 78.230 3322.425 78.560 3322.545 ;
        RECT 77.310 3322.255 78.560 3322.425 ;
        RECT 74.835 3321.795 75.850 3321.995 ;
        RECT 76.020 3321.615 76.430 3322.055 ;
        RECT 76.720 3321.825 76.970 3322.255 ;
        RECT 77.170 3321.615 77.490 3322.075 ;
        RECT 78.730 3322.005 78.900 3322.765 ;
        RECT 79.570 3322.705 79.900 3322.765 ;
        RECT 79.090 3322.535 79.420 3322.595 ;
        RECT 79.090 3322.265 79.750 3322.535 ;
        RECT 80.070 3322.210 80.260 3323.105 ;
        RECT 78.050 3321.835 78.900 3322.005 ;
        RECT 79.100 3321.615 79.760 3322.095 ;
        RECT 79.940 3321.880 80.260 3322.210 ;
        RECT 80.460 3322.855 80.710 3323.445 ;
        RECT 80.890 3323.365 81.175 3324.165 ;
        RECT 81.355 3323.185 81.610 3323.855 ;
        RECT 81.430 3322.890 81.610 3323.185 ;
        RECT 84.055 3323.235 84.225 3323.995 ;
        RECT 84.440 3323.405 84.770 3324.165 ;
        RECT 84.055 3323.065 84.770 3323.235 ;
        RECT 84.940 3323.090 85.195 3323.995 ;
        RECT 81.430 3322.885 83.980 3322.890 ;
        RECT 80.460 3322.525 81.260 3322.855 ;
        RECT 80.460 3321.875 80.710 3322.525 ;
        RECT 81.430 3322.515 84.320 3322.885 ;
        RECT 84.600 3322.855 84.770 3323.065 ;
        RECT 84.600 3322.525 84.855 3322.855 ;
        RECT 81.430 3322.490 83.980 3322.515 ;
        RECT 81.430 3322.325 81.610 3322.490 ;
        RECT 84.600 3322.335 84.770 3322.525 ;
        RECT 85.025 3322.360 85.195 3323.090 ;
        RECT 85.370 3323.990 88.180 3324.165 ;
        RECT 85.370 3323.015 85.630 3323.990 ;
        RECT 87.830 3323.540 88.180 3323.990 ;
        RECT 116.130 3323.070 116.530 3324.570 ;
        RECT 80.890 3321.615 81.175 3322.075 ;
        RECT 81.355 3321.795 81.610 3322.325 ;
        RECT 84.055 3322.165 84.770 3322.335 ;
        RECT 84.055 3321.785 84.225 3322.165 ;
        RECT 82.030 3321.615 83.880 3321.740 ;
        RECT 84.440 3321.615 84.770 3321.995 ;
        RECT 84.940 3321.785 85.195 3322.360 ;
        RECT 85.370 3321.615 85.630 3322.455 ;
        RECT 68.970 3321.445 85.720 3321.615 ;
        RECT 70.680 3321.290 72.430 3321.445 ;
        RECT 82.030 3321.290 83.880 3321.445 ;
        RECT 109.335 3320.770 109.505 3321.330 ;
        RECT 109.675 3320.985 110.225 3321.155 ;
        RECT 109.335 3320.440 109.885 3320.770 ;
        RECT 110.055 3320.610 110.225 3320.985 ;
        RECT 110.405 3320.890 110.775 3321.245 ;
        RECT 110.955 3320.985 111.885 3321.155 ;
        RECT 110.955 3320.610 111.125 3320.985 ;
        RECT 112.055 3320.770 112.225 3321.330 ;
        RECT 110.055 3320.440 111.125 3320.610 ;
        RECT 111.295 3320.440 112.225 3320.770 ;
        RECT 109.335 3319.840 109.505 3320.440 ;
        RECT 110.415 3320.355 110.745 3320.440 ;
        RECT 109.675 3320.185 110.250 3320.270 ;
        RECT 110.980 3320.185 111.885 3320.270 ;
        RECT 109.675 3320.015 111.885 3320.185 ;
        RECT 109.335 3319.580 110.345 3319.840 ;
        RECT 109.335 3319.490 109.505 3319.580 ;
        RECT 70.330 3319.125 77.480 3319.140 ;
        RECT 69.120 3318.955 77.480 3319.125 ;
        RECT 68.430 3318.340 68.830 3318.840 ;
        RECT 69.245 3317.815 69.475 3318.955 ;
        RECT 70.145 3318.790 77.480 3318.955 ;
        RECT 69.645 3317.805 69.975 3318.785 ;
        RECT 70.145 3317.815 70.355 3318.790 ;
        RECT 77.130 3318.655 77.480 3318.790 ;
        RECT 77.130 3318.485 80.350 3318.655 ;
        RECT 81.710 3318.640 83.550 3318.655 ;
        RECT 87.830 3318.640 88.180 3319.090 ;
        RECT 109.680 3318.770 110.180 3319.170 ;
        RECT 81.710 3318.485 88.180 3318.640 ;
        RECT 64.180 3317.320 68.880 3317.720 ;
        RECT 69.225 3317.395 69.555 3317.645 ;
        RECT 69.725 3317.590 69.975 3317.805 ;
        RECT 77.215 3317.635 77.595 3318.315 ;
        RECT 78.185 3317.635 78.355 3318.485 ;
        RECT 78.525 3317.805 78.855 3318.315 ;
        RECT 79.025 3317.975 79.195 3318.485 ;
        RECT 79.365 3317.805 79.765 3318.315 ;
        RECT 78.525 3317.635 79.765 3317.805 ;
        RECT 69.725 3317.420 69.980 3317.590 ;
        RECT 68.430 3316.590 68.830 3317.090 ;
        RECT 69.245 3316.405 69.475 3317.225 ;
        RECT 69.725 3317.205 69.975 3317.420 ;
        RECT 69.645 3316.575 69.975 3317.205 ;
        RECT 70.145 3316.590 70.355 3317.225 ;
        RECT 77.215 3316.675 77.385 3317.635 ;
        RECT 77.555 3317.295 78.860 3317.465 ;
        RECT 79.945 3317.385 80.265 3318.315 ;
        RECT 80.880 3317.590 81.280 3318.090 ;
        RECT 81.885 3317.555 82.055 3318.315 ;
        RECT 82.270 3317.725 82.600 3318.485 ;
        RECT 81.885 3317.385 82.600 3317.555 ;
        RECT 82.770 3317.410 83.025 3318.315 ;
        RECT 77.555 3316.845 77.800 3317.295 ;
        RECT 77.970 3316.925 78.520 3317.125 ;
        RECT 78.690 3317.095 78.860 3317.295 ;
        RECT 79.635 3317.240 80.265 3317.385 ;
        RECT 79.635 3317.190 81.480 3317.240 ;
        RECT 81.795 3317.190 82.150 3317.205 ;
        RECT 78.690 3316.925 79.065 3317.095 ;
        RECT 79.235 3316.675 79.465 3317.175 ;
        RECT 70.145 3316.405 75.030 3316.590 ;
        RECT 77.215 3316.505 79.465 3316.675 ;
        RECT 79.635 3316.990 82.150 3317.190 ;
        RECT 69.120 3316.240 75.030 3316.405 ;
        RECT 69.120 3316.235 70.500 3316.240 ;
        RECT 74.680 3316.040 75.030 3316.240 ;
        RECT 77.265 3316.040 77.595 3316.325 ;
        RECT 77.765 3316.185 77.935 3316.505 ;
        RECT 79.635 3316.335 79.805 3316.990 ;
        RECT 81.795 3316.835 82.150 3316.990 ;
        RECT 82.430 3317.175 82.600 3317.385 ;
        RECT 82.430 3316.845 82.685 3317.175 ;
        RECT 74.680 3315.935 77.595 3316.040 ;
        RECT 78.105 3315.935 78.435 3316.325 ;
        RECT 78.850 3316.165 79.805 3316.335 ;
        RECT 79.975 3315.935 80.265 3316.770 ;
        RECT 82.430 3316.655 82.600 3316.845 ;
        RECT 82.855 3316.680 83.025 3317.410 ;
        RECT 83.200 3318.290 88.180 3318.485 ;
        RECT 83.200 3317.335 83.460 3318.290 ;
        RECT 87.830 3317.890 88.180 3318.290 ;
        RECT 110.530 3318.670 110.730 3320.015 ;
        RECT 112.055 3319.840 112.225 3320.440 ;
        RECT 110.905 3319.580 112.225 3319.840 ;
        RECT 112.055 3319.490 112.225 3319.580 ;
        RECT 116.830 3319.520 117.230 3323.520 ;
        RECT 111.080 3318.870 111.580 3319.270 ;
        RECT 117.230 3319.070 117.530 3319.120 ;
        RECT 112.930 3318.670 117.530 3319.070 ;
        RECT 110.530 3318.270 113.330 3318.670 ;
        RECT 117.230 3318.620 117.530 3318.670 ;
        RECT 109.335 3317.905 109.505 3318.030 ;
        RECT 110.530 3317.925 110.730 3318.270 ;
        RECT 109.335 3317.675 110.325 3317.905 ;
        RECT 84.480 3316.870 90.030 3317.270 ;
        RECT 109.335 3317.005 109.505 3317.675 ;
        RECT 110.495 3317.595 110.745 3317.925 ;
        RECT 112.055 3317.905 112.225 3318.030 ;
        RECT 110.915 3317.675 112.225 3317.905 ;
        RECT 109.675 3317.425 110.305 3317.505 ;
        RECT 110.905 3317.425 111.885 3317.505 ;
        RECT 109.675 3317.175 111.885 3317.425 ;
        RECT 112.055 3317.005 112.225 3317.675 ;
        RECT 117.730 3317.920 118.130 3323.520 ;
        RECT 118.630 3319.520 119.030 3324.570 ;
        RECT 120.930 3322.920 121.330 3323.420 ;
        RECT 118.330 3318.620 118.630 3319.120 ;
        RECT 121.630 3317.920 122.030 3323.370 ;
        RECT 122.530 3321.370 122.930 3325.570 ;
        RECT 123.430 3321.370 123.830 3323.370 ;
        RECT 125.480 3321.370 125.880 3323.370 ;
        RECT 126.380 3321.370 126.780 3325.570 ;
        RECT 129.980 3325.070 130.380 3325.570 ;
        RECT 129.980 3324.570 131.080 3325.070 ;
        RECT 122.230 3320.470 123.230 3320.970 ;
        RECT 126.180 3320.470 127.030 3320.970 ;
        RECT 117.730 3317.520 122.030 3317.920 ;
        RECT 122.530 3317.120 122.930 3320.470 ;
        RECT 127.280 3318.270 127.680 3323.370 ;
        RECT 129.980 3322.920 130.380 3324.570 ;
        RECT 127.980 3321.320 128.380 3321.820 ;
        RECT 130.680 3319.470 131.080 3324.570 ;
        RECT 131.080 3318.570 131.380 3319.070 ;
        RECT 131.580 3318.270 131.980 3323.470 ;
        RECT 132.480 3319.470 132.880 3323.470 ;
        RECT 132.180 3318.570 132.480 3319.070 ;
        RECT 134.080 3318.270 134.580 3328.720 ;
        RECT 148.580 3328.745 149.605 3328.995 ;
        RECT 139.980 3327.720 140.480 3328.320 ;
        RECT 146.530 3328.165 148.180 3328.320 ;
        RECT 143.770 3327.995 148.180 3328.165 ;
        RECT 139.980 3327.220 141.080 3327.720 ;
        RECT 143.030 3327.220 143.430 3327.720 ;
        RECT 139.980 3320.270 140.480 3327.220 ;
        RECT 143.865 3327.015 144.195 3327.825 ;
        RECT 144.365 3327.195 144.605 3327.995 ;
        RECT 143.865 3326.845 144.580 3327.015 ;
        RECT 143.860 3326.670 144.240 3326.675 ;
        RECT 142.280 3326.470 144.240 3326.670 ;
        RECT 142.280 3324.320 142.580 3326.470 ;
        RECT 143.860 3326.435 144.240 3326.470 ;
        RECT 144.410 3326.605 144.580 3326.845 ;
        RECT 144.785 3326.975 144.955 3327.825 ;
        RECT 145.125 3327.195 145.455 3327.995 ;
        RECT 145.625 3326.975 145.795 3327.825 ;
        RECT 144.785 3326.805 145.795 3326.975 ;
        RECT 145.965 3326.845 146.295 3327.995 ;
        RECT 146.530 3327.870 148.180 3327.995 ;
        RECT 148.580 3327.470 148.830 3328.745 ;
        RECT 158.830 3328.420 159.230 3332.170 ;
        RECT 149.170 3327.995 158.830 3328.165 ;
        RECT 146.530 3327.220 148.830 3327.470 ;
        RECT 149.345 3327.325 149.515 3327.825 ;
        RECT 149.685 3327.495 150.015 3327.995 ;
        RECT 145.300 3326.670 145.795 3326.805 ;
        RECT 146.530 3326.670 146.805 3327.220 ;
        RECT 149.345 3327.155 150.010 3327.325 ;
        RECT 144.410 3326.435 144.910 3326.605 ;
        RECT 144.410 3326.265 144.580 3326.435 ;
        RECT 145.300 3326.420 146.805 3326.670 ;
        RECT 145.300 3326.265 145.795 3326.420 ;
        RECT 149.260 3326.335 149.610 3326.985 ;
        RECT 143.945 3326.095 144.580 3326.265 ;
        RECT 144.785 3326.095 145.795 3326.265 ;
        RECT 143.030 3325.420 143.430 3325.920 ;
        RECT 143.945 3325.615 144.115 3326.095 ;
        RECT 144.295 3325.445 144.535 3325.925 ;
        RECT 144.785 3325.615 144.955 3326.095 ;
        RECT 145.125 3325.445 145.455 3325.925 ;
        RECT 145.625 3325.615 145.795 3326.095 ;
        RECT 145.965 3325.445 146.295 3326.245 ;
        RECT 149.780 3326.165 150.010 3327.155 ;
        RECT 149.345 3325.995 150.010 3326.165 ;
        RECT 149.345 3325.705 149.515 3325.995 ;
        RECT 146.530 3325.445 149.180 3325.620 ;
        RECT 149.685 3325.445 150.015 3325.825 ;
        RECT 150.185 3325.705 150.370 3327.825 ;
        RECT 150.610 3327.535 150.875 3327.995 ;
        RECT 151.045 3327.400 151.295 3327.825 ;
        RECT 151.505 3327.550 152.610 3327.720 ;
        RECT 150.990 3327.270 151.295 3327.400 ;
        RECT 150.540 3326.075 150.820 3327.025 ;
        RECT 150.990 3326.165 151.160 3327.270 ;
        RECT 151.330 3326.485 151.570 3327.080 ;
        RECT 151.740 3327.015 152.270 3327.380 ;
        RECT 151.740 3326.315 151.910 3327.015 ;
        RECT 152.440 3326.935 152.610 3327.550 ;
        RECT 152.780 3327.195 152.950 3327.995 ;
        RECT 153.120 3327.495 153.370 3327.825 ;
        RECT 153.595 3327.525 154.480 3327.695 ;
        RECT 152.440 3326.845 152.950 3326.935 ;
        RECT 150.990 3326.035 151.215 3326.165 ;
        RECT 151.385 3326.095 151.910 3326.315 ;
        RECT 152.080 3326.675 152.950 3326.845 ;
        RECT 150.625 3325.445 150.875 3325.905 ;
        RECT 151.045 3325.895 151.215 3326.035 ;
        RECT 152.080 3325.895 152.250 3326.675 ;
        RECT 152.780 3326.605 152.950 3326.675 ;
        RECT 152.460 3326.425 152.660 3326.455 ;
        RECT 153.120 3326.425 153.290 3327.495 ;
        RECT 153.460 3326.605 153.650 3327.325 ;
        RECT 152.460 3326.125 153.290 3326.425 ;
        RECT 153.820 3326.395 154.140 3327.355 ;
        RECT 151.045 3325.725 151.380 3325.895 ;
        RECT 151.575 3325.725 152.250 3325.895 ;
        RECT 152.570 3325.445 152.940 3325.945 ;
        RECT 153.120 3325.895 153.290 3326.125 ;
        RECT 153.675 3326.065 154.140 3326.395 ;
        RECT 154.310 3326.685 154.480 3327.525 ;
        RECT 154.660 3327.495 154.975 3327.995 ;
        RECT 155.210 3327.265 155.550 3327.825 ;
        RECT 154.650 3326.890 155.550 3327.265 ;
        RECT 155.720 3326.985 155.890 3327.995 ;
        RECT 155.360 3326.685 155.550 3326.890 ;
        RECT 156.060 3326.935 156.390 3327.780 ;
        RECT 156.560 3327.080 156.735 3327.995 ;
        RECT 157.075 3327.075 157.405 3327.805 ;
        RECT 156.060 3326.855 156.470 3326.935 ;
        RECT 156.235 3326.805 156.470 3326.855 ;
        RECT 154.310 3326.355 155.190 3326.685 ;
        RECT 155.360 3326.355 156.110 3326.685 ;
        RECT 154.310 3325.895 154.480 3326.355 ;
        RECT 155.360 3326.185 155.560 3326.355 ;
        RECT 156.280 3326.225 156.470 3326.805 ;
        RECT 156.225 3326.185 156.470 3326.225 ;
        RECT 153.120 3325.725 153.525 3325.895 ;
        RECT 153.695 3325.725 154.480 3325.895 ;
        RECT 154.755 3325.445 154.965 3325.975 ;
        RECT 155.230 3325.660 155.560 3326.185 ;
        RECT 156.070 3326.100 156.470 3326.185 ;
        RECT 157.135 3326.685 157.405 3327.075 ;
        RECT 157.595 3326.855 157.810 3327.995 ;
        RECT 157.980 3326.855 158.315 3327.825 ;
        RECT 158.485 3326.855 158.735 3327.995 ;
        RECT 159.180 3326.870 159.680 3327.270 ;
        RECT 157.135 3326.355 157.930 3326.685 ;
        RECT 158.100 3326.670 158.315 3326.855 ;
        RECT 158.100 3326.470 160.280 3326.670 ;
        RECT 155.730 3325.445 155.900 3326.055 ;
        RECT 156.070 3325.665 156.400 3326.100 ;
        RECT 157.135 3325.975 157.335 3326.355 ;
        RECT 158.100 3326.245 158.315 3326.470 ;
        RECT 158.930 3326.320 160.280 3326.470 ;
        RECT 156.570 3325.445 156.740 3325.960 ;
        RECT 157.075 3325.705 157.335 3325.975 ;
        RECT 157.560 3325.445 157.890 3326.185 ;
        RECT 158.060 3325.625 158.315 3326.245 ;
        RECT 158.485 3325.445 158.735 3326.265 ;
        RECT 159.080 3325.720 159.580 3326.120 ;
        RECT 143.770 3325.275 158.830 3325.445 ;
        RECT 146.530 3325.120 149.180 3325.275 ;
        RECT 159.880 3324.320 160.280 3326.320 ;
        RECT 142.280 3323.920 160.280 3324.320 ;
        RECT 157.880 3320.665 159.230 3320.820 ;
        RECT 145.970 3320.495 148.270 3320.665 ;
        RECT 150.570 3320.495 159.230 3320.665 ;
        RECT 139.980 3319.770 141.080 3320.270 ;
        RECT 144.030 3319.770 144.430 3320.270 ;
        RECT 139.980 3319.170 140.480 3319.770 ;
        RECT 146.100 3319.355 146.365 3320.495 ;
        RECT 146.535 3319.525 146.865 3320.325 ;
        RECT 147.035 3319.695 147.205 3320.495 ;
        RECT 147.375 3319.545 147.705 3320.325 ;
        RECT 147.875 3320.035 148.085 3320.495 ;
        RECT 150.745 3319.825 150.915 3320.325 ;
        RECT 151.085 3319.995 151.415 3320.495 ;
        RECT 150.745 3319.655 151.410 3319.825 ;
        RECT 147.375 3319.525 148.140 3319.545 ;
        RECT 146.535 3319.470 148.140 3319.525 ;
        RECT 150.660 3319.470 151.010 3319.485 ;
        RECT 146.535 3319.355 151.010 3319.470 ;
        RECT 127.280 3317.770 134.580 3318.270 ;
        RECT 137.830 3318.620 138.330 3318.970 ;
        RECT 146.075 3318.935 147.705 3319.185 ;
        RECT 147.875 3319.070 151.010 3319.355 ;
        RECT 147.875 3318.765 148.140 3319.070 ;
        RECT 150.660 3318.835 151.010 3319.070 ;
        RECT 137.830 3318.120 144.430 3318.620 ;
        RECT 146.535 3318.585 148.140 3318.765 ;
        RECT 151.180 3318.665 151.410 3319.655 ;
        RECT 137.830 3317.770 138.330 3318.120 ;
        RECT 146.100 3317.945 146.365 3318.405 ;
        RECT 146.535 3318.115 146.865 3318.585 ;
        RECT 147.035 3317.945 147.205 3318.405 ;
        RECT 147.375 3318.115 147.705 3318.585 ;
        RECT 147.875 3317.945 148.125 3318.410 ;
        RECT 149.180 3318.170 149.730 3318.620 ;
        RECT 150.745 3318.495 151.410 3318.665 ;
        RECT 150.745 3318.205 150.915 3318.495 ;
        RECT 145.970 3317.775 148.270 3317.945 ;
        RECT 149.355 3317.295 149.605 3318.170 ;
        RECT 151.085 3317.945 151.415 3318.325 ;
        RECT 151.585 3318.205 151.770 3320.325 ;
        RECT 152.010 3320.035 152.275 3320.495 ;
        RECT 152.445 3319.900 152.695 3320.325 ;
        RECT 152.905 3320.050 154.010 3320.220 ;
        RECT 152.390 3319.770 152.695 3319.900 ;
        RECT 151.940 3318.575 152.220 3319.525 ;
        RECT 152.390 3318.665 152.560 3319.770 ;
        RECT 152.730 3318.985 152.970 3319.580 ;
        RECT 153.140 3319.515 153.670 3319.880 ;
        RECT 153.140 3318.815 153.310 3319.515 ;
        RECT 153.840 3319.435 154.010 3320.050 ;
        RECT 154.180 3319.695 154.350 3320.495 ;
        RECT 154.520 3319.995 154.770 3320.325 ;
        RECT 154.995 3320.025 155.880 3320.195 ;
        RECT 153.840 3319.345 154.350 3319.435 ;
        RECT 152.390 3318.535 152.615 3318.665 ;
        RECT 152.785 3318.595 153.310 3318.815 ;
        RECT 153.480 3319.175 154.350 3319.345 ;
        RECT 152.025 3317.945 152.275 3318.405 ;
        RECT 152.445 3318.395 152.615 3318.535 ;
        RECT 153.480 3318.395 153.650 3319.175 ;
        RECT 154.180 3319.105 154.350 3319.175 ;
        RECT 153.860 3318.925 154.060 3318.955 ;
        RECT 154.520 3318.925 154.690 3319.995 ;
        RECT 154.860 3319.105 155.050 3319.825 ;
        RECT 153.860 3318.625 154.690 3318.925 ;
        RECT 155.220 3318.895 155.540 3319.855 ;
        RECT 152.445 3318.225 152.780 3318.395 ;
        RECT 152.975 3318.225 153.650 3318.395 ;
        RECT 153.970 3317.945 154.340 3318.445 ;
        RECT 154.520 3318.395 154.690 3318.625 ;
        RECT 155.075 3318.565 155.540 3318.895 ;
        RECT 155.710 3319.185 155.880 3320.025 ;
        RECT 156.060 3319.995 156.375 3320.495 ;
        RECT 156.605 3319.765 156.945 3320.325 ;
        RECT 156.050 3319.390 156.945 3319.765 ;
        RECT 157.115 3319.485 157.285 3320.495 ;
        RECT 157.880 3320.470 159.230 3320.495 ;
        RECT 156.755 3319.185 156.945 3319.390 ;
        RECT 157.455 3319.435 157.785 3320.280 ;
        RECT 157.455 3319.355 157.845 3319.435 ;
        RECT 157.630 3319.305 157.845 3319.355 ;
        RECT 155.710 3318.855 156.585 3319.185 ;
        RECT 156.755 3318.855 157.505 3319.185 ;
        RECT 155.710 3318.395 155.880 3318.855 ;
        RECT 156.755 3318.685 156.955 3318.855 ;
        RECT 157.675 3318.725 157.845 3319.305 ;
        RECT 157.620 3318.685 157.845 3318.725 ;
        RECT 154.520 3318.225 154.925 3318.395 ;
        RECT 155.095 3318.225 155.880 3318.395 ;
        RECT 156.155 3317.945 156.365 3318.475 ;
        RECT 156.625 3318.160 156.955 3318.685 ;
        RECT 157.465 3318.600 157.845 3318.685 ;
        RECT 157.125 3317.945 157.295 3318.555 ;
        RECT 157.465 3318.165 157.795 3318.600 ;
        RECT 150.570 3317.775 157.930 3317.945 ;
        RECT 109.335 3316.795 110.325 3317.005 ;
        RECT 110.915 3316.795 112.225 3317.005 ;
        RECT 80.780 3316.090 81.280 3316.490 ;
        RECT 81.885 3316.485 82.600 3316.655 ;
        RECT 81.885 3316.105 82.055 3316.485 ;
        RECT 82.270 3315.935 82.600 3316.315 ;
        RECT 82.770 3316.105 83.025 3316.680 ;
        RECT 83.200 3315.935 83.460 3316.775 ;
        RECT 109.335 3316.650 109.505 3316.795 ;
        RECT 112.055 3316.650 112.225 3316.795 ;
        RECT 112.930 3316.620 132.880 3317.120 ;
        RECT 148.580 3317.045 149.605 3317.295 ;
        RECT 112.930 3316.020 113.430 3316.620 ;
        RECT 146.530 3316.465 148.180 3316.620 ;
        RECT 143.770 3316.295 148.180 3316.465 ;
        RECT 74.680 3315.765 80.350 3315.935 ;
        RECT 81.710 3315.765 83.550 3315.935 ;
        RECT 74.680 3315.690 77.330 3315.765 ;
        RECT 71.230 3313.965 72.530 3314.090 ;
        RECT 74.680 3313.965 75.030 3315.690 ;
        RECT 110.780 3315.520 113.430 3316.020 ;
        RECT 116.480 3315.470 121.330 3315.870 ;
        RECT 143.030 3315.520 143.430 3316.020 ;
        RECT 143.865 3315.315 144.195 3316.125 ;
        RECT 144.365 3315.495 144.605 3316.295 ;
        RECT 143.865 3315.145 144.580 3315.315 ;
        RECT 143.860 3314.970 144.240 3314.975 ;
        RECT 118.360 3314.630 132.380 3314.800 ;
        RECT 82.080 3313.965 84.230 3313.990 ;
        RECT 69.980 3313.795 85.880 3313.965 ;
        RECT 70.125 3312.975 70.335 3313.795 ;
        RECT 71.005 3313.640 72.530 3313.795 ;
        RECT 70.505 3312.995 70.835 3313.625 ;
        RECT 70.505 3312.395 70.755 3312.995 ;
        RECT 71.005 3312.975 71.235 3313.640 ;
        RECT 72.910 3313.085 73.165 3313.615 ;
        RECT 73.345 3313.335 73.630 3313.795 ;
        RECT 70.925 3312.800 71.255 3312.805 ;
        RECT 72.910 3312.800 73.090 3313.085 ;
        RECT 73.810 3312.885 74.060 3313.535 ;
        RECT 70.925 3312.560 73.090 3312.800 ;
        RECT 70.925 3312.555 71.255 3312.560 ;
        RECT 70.125 3311.245 70.335 3312.385 ;
        RECT 70.505 3311.415 70.835 3312.395 ;
        RECT 71.005 3311.245 71.235 3312.385 ;
        RECT 72.910 3312.225 73.090 3312.560 ;
        RECT 73.260 3312.555 74.060 3312.885 ;
        RECT 71.830 3311.640 72.230 3312.140 ;
        RECT 72.910 3311.555 73.165 3312.225 ;
        RECT 73.345 3311.245 73.630 3312.045 ;
        RECT 73.810 3311.965 74.060 3312.555 ;
        RECT 74.260 3313.200 74.580 3313.530 ;
        RECT 74.760 3313.315 75.420 3313.795 ;
        RECT 75.620 3313.405 76.470 3313.575 ;
        RECT 74.260 3312.305 74.450 3313.200 ;
        RECT 74.770 3312.875 75.430 3313.145 ;
        RECT 75.100 3312.815 75.430 3312.875 ;
        RECT 74.620 3312.645 74.950 3312.705 ;
        RECT 75.620 3312.645 75.790 3313.405 ;
        RECT 77.030 3313.335 77.350 3313.795 ;
        RECT 77.550 3313.155 77.800 3313.585 ;
        RECT 78.090 3313.355 78.500 3313.795 ;
        RECT 78.670 3313.415 79.685 3313.615 ;
        RECT 75.960 3312.985 77.210 3313.155 ;
        RECT 75.960 3312.865 76.290 3312.985 ;
        RECT 74.620 3312.475 76.520 3312.645 ;
        RECT 74.260 3312.135 76.180 3312.305 ;
        RECT 74.260 3312.115 74.580 3312.135 ;
        RECT 73.810 3311.455 74.140 3311.965 ;
        RECT 74.410 3311.505 74.580 3312.115 ;
        RECT 76.350 3311.965 76.520 3312.475 ;
        RECT 76.690 3312.405 76.870 3312.815 ;
        RECT 77.040 3312.225 77.210 3312.985 ;
        RECT 74.750 3311.245 75.080 3311.935 ;
        RECT 75.310 3311.795 76.520 3311.965 ;
        RECT 76.690 3311.915 77.210 3312.225 ;
        RECT 77.380 3312.815 77.800 3313.155 ;
        RECT 78.090 3312.815 78.500 3313.145 ;
        RECT 77.380 3312.045 77.570 3312.815 ;
        RECT 78.670 3312.685 78.840 3313.415 ;
        RECT 79.985 3313.245 80.155 3313.575 ;
        RECT 80.325 3313.415 80.655 3313.795 ;
        RECT 79.010 3312.865 79.360 3313.235 ;
        RECT 78.670 3312.645 79.090 3312.685 ;
        RECT 77.740 3312.475 79.090 3312.645 ;
        RECT 77.740 3312.315 77.990 3312.475 ;
        RECT 78.500 3312.045 78.750 3312.305 ;
        RECT 77.380 3311.795 78.750 3312.045 ;
        RECT 75.310 3311.505 75.550 3311.795 ;
        RECT 76.350 3311.715 76.520 3311.795 ;
        RECT 75.750 3311.245 76.170 3311.625 ;
        RECT 76.350 3311.465 76.980 3311.715 ;
        RECT 77.450 3311.245 77.780 3311.625 ;
        RECT 77.950 3311.505 78.120 3311.795 ;
        RECT 78.920 3311.630 79.090 3312.475 ;
        RECT 79.540 3312.305 79.760 3313.175 ;
        RECT 79.985 3313.055 80.680 3313.245 ;
        RECT 79.260 3311.925 79.760 3312.305 ;
        RECT 79.930 3312.255 80.340 3312.875 ;
        RECT 80.510 3312.085 80.680 3313.055 ;
        RECT 79.985 3311.915 80.680 3312.085 ;
        RECT 78.300 3311.245 78.680 3311.625 ;
        RECT 78.920 3311.460 79.750 3311.630 ;
        RECT 79.985 3311.415 80.155 3311.915 ;
        RECT 80.325 3311.245 80.655 3311.745 ;
        RECT 80.870 3311.415 81.095 3313.535 ;
        RECT 81.265 3313.415 81.595 3313.795 ;
        RECT 82.080 3313.640 84.390 3313.795 ;
        RECT 81.765 3313.245 81.935 3313.535 ;
        RECT 81.270 3313.075 81.935 3313.245 ;
        RECT 83.180 3313.240 83.680 3313.640 ;
        RECT 81.270 3312.085 81.500 3313.075 ;
        RECT 84.130 3312.955 84.390 3313.640 ;
        RECT 84.565 3313.050 84.820 3313.625 ;
        RECT 84.990 3313.415 85.320 3313.795 ;
        RECT 85.535 3313.245 85.705 3313.625 ;
        RECT 84.990 3313.075 85.705 3313.245 ;
        RECT 81.670 3312.890 82.020 3312.905 ;
        RECT 81.670 3312.540 83.580 3312.890 ;
        RECT 81.670 3312.255 82.020 3312.540 ;
        RECT 81.270 3311.915 81.935 3312.085 ;
        RECT 81.265 3311.245 81.595 3311.745 ;
        RECT 81.765 3311.415 81.935 3311.915 ;
        RECT 84.130 3311.245 84.390 3312.395 ;
        RECT 84.565 3312.320 84.735 3313.050 ;
        RECT 84.990 3312.885 85.160 3313.075 ;
        RECT 98.180 3313.070 98.780 3313.670 ;
        RECT 118.360 3313.470 118.530 3314.630 ;
        RECT 131.630 3314.150 131.930 3314.170 ;
        RECT 119.010 3313.800 121.170 3314.150 ;
        RECT 129.570 3313.800 131.930 3314.150 ;
        RECT 118.280 3313.320 118.680 3313.470 ;
        RECT 131.630 3313.320 131.930 3313.800 ;
        RECT 132.210 3313.320 132.380 3314.630 ;
        RECT 118.280 3313.150 132.380 3313.320 ;
        RECT 142.280 3314.770 144.240 3314.970 ;
        RECT 118.280 3313.070 118.680 3313.150 ;
        RECT 86.080 3312.900 98.780 3313.070 ;
        RECT 84.905 3312.555 85.160 3312.885 ;
        RECT 84.990 3312.345 85.160 3312.555 ;
        RECT 85.440 3312.520 98.780 3312.900 ;
        RECT 86.080 3312.470 98.780 3312.520 ;
        RECT 142.280 3312.620 142.580 3314.770 ;
        RECT 143.860 3314.735 144.240 3314.770 ;
        RECT 144.410 3314.905 144.580 3315.145 ;
        RECT 144.785 3315.275 144.955 3316.125 ;
        RECT 145.125 3315.495 145.455 3316.295 ;
        RECT 145.625 3315.275 145.795 3316.125 ;
        RECT 144.785 3315.105 145.795 3315.275 ;
        RECT 145.965 3315.145 146.295 3316.295 ;
        RECT 146.530 3316.170 148.180 3316.295 ;
        RECT 148.580 3315.770 148.830 3317.045 ;
        RECT 158.830 3316.720 159.230 3320.470 ;
        RECT 159.580 3316.770 164.030 3317.270 ;
        RECT 149.170 3316.295 158.830 3316.465 ;
        RECT 159.580 3316.370 160.080 3316.770 ;
        RECT 146.530 3315.520 148.830 3315.770 ;
        RECT 149.345 3315.625 149.515 3316.125 ;
        RECT 149.685 3315.795 150.015 3316.295 ;
        RECT 145.300 3314.970 145.795 3315.105 ;
        RECT 146.530 3314.970 146.805 3315.520 ;
        RECT 149.345 3315.455 150.010 3315.625 ;
        RECT 144.410 3314.735 144.910 3314.905 ;
        RECT 144.410 3314.565 144.580 3314.735 ;
        RECT 145.300 3314.720 146.805 3314.970 ;
        RECT 145.300 3314.565 145.795 3314.720 ;
        RECT 149.260 3314.635 149.610 3315.285 ;
        RECT 143.945 3314.395 144.580 3314.565 ;
        RECT 144.785 3314.395 145.795 3314.565 ;
        RECT 143.030 3313.720 143.430 3314.220 ;
        RECT 143.945 3313.915 144.115 3314.395 ;
        RECT 144.295 3313.745 144.535 3314.225 ;
        RECT 144.785 3313.915 144.955 3314.395 ;
        RECT 145.125 3313.745 145.455 3314.225 ;
        RECT 145.625 3313.915 145.795 3314.395 ;
        RECT 145.965 3313.745 146.295 3314.545 ;
        RECT 149.780 3314.465 150.010 3315.455 ;
        RECT 149.345 3314.295 150.010 3314.465 ;
        RECT 149.345 3314.005 149.515 3314.295 ;
        RECT 146.530 3313.745 149.180 3313.920 ;
        RECT 149.685 3313.745 150.015 3314.125 ;
        RECT 150.185 3314.005 150.370 3316.125 ;
        RECT 150.610 3315.835 150.875 3316.295 ;
        RECT 151.045 3315.700 151.295 3316.125 ;
        RECT 151.505 3315.850 152.610 3316.020 ;
        RECT 150.990 3315.570 151.295 3315.700 ;
        RECT 150.540 3314.375 150.820 3315.325 ;
        RECT 150.990 3314.465 151.160 3315.570 ;
        RECT 151.330 3314.785 151.570 3315.380 ;
        RECT 151.740 3315.315 152.270 3315.680 ;
        RECT 151.740 3314.615 151.910 3315.315 ;
        RECT 152.440 3315.235 152.610 3315.850 ;
        RECT 152.780 3315.495 152.950 3316.295 ;
        RECT 153.120 3315.795 153.370 3316.125 ;
        RECT 153.595 3315.825 154.480 3315.995 ;
        RECT 152.440 3315.145 152.950 3315.235 ;
        RECT 150.990 3314.335 151.215 3314.465 ;
        RECT 151.385 3314.395 151.910 3314.615 ;
        RECT 152.080 3314.975 152.950 3315.145 ;
        RECT 150.625 3313.745 150.875 3314.205 ;
        RECT 151.045 3314.195 151.215 3314.335 ;
        RECT 152.080 3314.195 152.250 3314.975 ;
        RECT 152.780 3314.905 152.950 3314.975 ;
        RECT 152.460 3314.725 152.660 3314.755 ;
        RECT 153.120 3314.725 153.290 3315.795 ;
        RECT 153.460 3314.905 153.650 3315.625 ;
        RECT 152.460 3314.425 153.290 3314.725 ;
        RECT 153.820 3314.695 154.140 3315.655 ;
        RECT 151.045 3314.025 151.380 3314.195 ;
        RECT 151.575 3314.025 152.250 3314.195 ;
        RECT 152.570 3313.745 152.940 3314.245 ;
        RECT 153.120 3314.195 153.290 3314.425 ;
        RECT 153.675 3314.365 154.140 3314.695 ;
        RECT 154.310 3314.985 154.480 3315.825 ;
        RECT 154.660 3315.795 154.975 3316.295 ;
        RECT 155.210 3315.565 155.550 3316.125 ;
        RECT 154.650 3315.190 155.550 3315.565 ;
        RECT 155.720 3315.285 155.890 3316.295 ;
        RECT 155.360 3314.985 155.550 3315.190 ;
        RECT 156.060 3315.235 156.390 3316.080 ;
        RECT 156.560 3315.380 156.735 3316.295 ;
        RECT 157.075 3315.375 157.405 3316.105 ;
        RECT 156.060 3315.155 156.470 3315.235 ;
        RECT 156.235 3315.105 156.470 3315.155 ;
        RECT 154.310 3314.655 155.190 3314.985 ;
        RECT 155.360 3314.655 156.110 3314.985 ;
        RECT 154.310 3314.195 154.480 3314.655 ;
        RECT 155.360 3314.485 155.560 3314.655 ;
        RECT 156.280 3314.525 156.470 3315.105 ;
        RECT 156.225 3314.485 156.470 3314.525 ;
        RECT 153.120 3314.025 153.525 3314.195 ;
        RECT 153.695 3314.025 154.480 3314.195 ;
        RECT 154.755 3313.745 154.965 3314.275 ;
        RECT 155.230 3313.960 155.560 3314.485 ;
        RECT 156.070 3314.400 156.470 3314.485 ;
        RECT 157.135 3314.985 157.405 3315.375 ;
        RECT 157.595 3315.155 157.810 3316.295 ;
        RECT 157.980 3315.155 158.315 3316.125 ;
        RECT 158.485 3315.155 158.735 3316.295 ;
        RECT 159.180 3315.170 159.680 3315.570 ;
        RECT 157.135 3314.655 157.930 3314.985 ;
        RECT 158.100 3314.970 158.315 3315.155 ;
        RECT 158.100 3314.770 160.280 3314.970 ;
        RECT 155.730 3313.745 155.900 3314.355 ;
        RECT 156.070 3313.965 156.400 3314.400 ;
        RECT 157.135 3314.275 157.335 3314.655 ;
        RECT 158.100 3314.545 158.315 3314.770 ;
        RECT 158.930 3314.620 160.280 3314.770 ;
        RECT 156.570 3313.745 156.740 3314.260 ;
        RECT 157.075 3314.005 157.335 3314.275 ;
        RECT 157.560 3313.745 157.890 3314.485 ;
        RECT 158.060 3313.925 158.315 3314.545 ;
        RECT 158.485 3313.745 158.735 3314.565 ;
        RECT 159.080 3314.020 159.580 3314.420 ;
        RECT 143.770 3313.575 158.830 3313.745 ;
        RECT 146.530 3313.420 149.180 3313.575 ;
        RECT 159.880 3312.620 160.280 3314.620 ;
        RECT 84.565 3311.415 84.820 3312.320 ;
        RECT 84.990 3312.175 85.705 3312.345 ;
        RECT 142.280 3312.220 160.280 3312.620 ;
        RECT 84.990 3311.245 85.320 3312.005 ;
        RECT 85.535 3311.415 85.705 3312.175 ;
        RECT 87.830 3311.290 88.180 3311.740 ;
        RECT 85.830 3311.245 88.180 3311.290 ;
        RECT 69.980 3311.075 71.360 3311.245 ;
        RECT 72.450 3311.075 82.110 3311.245 ;
        RECT 84.040 3311.075 88.180 3311.245 ;
        RECT 69.980 3310.920 71.280 3311.075 ;
        RECT 85.830 3310.940 88.180 3311.075 ;
        RECT 66.180 3309.720 71.280 3310.920 ;
        RECT 68.980 3308.820 71.280 3309.720 ;
        RECT 163.530 3306.520 164.030 3316.770 ;
        RECT 163.180 3306.120 164.030 3306.520 ;
      LAYER met1 ;
        RECT 74.630 3396.570 76.630 3396.970 ;
        RECT 94.280 3396.570 96.280 3396.970 ;
        RECT 133.380 3396.570 135.380 3396.970 ;
        RECT 157.530 3396.570 159.530 3396.970 ;
        RECT 71.280 3395.220 71.680 3395.720 ;
        RECT 80.780 3395.220 81.180 3395.720 ;
        RECT 86.230 3395.220 86.630 3395.720 ;
        RECT 91.680 3395.220 92.080 3395.720 ;
        RECT 101.280 3395.220 101.680 3395.720 ;
        RECT 110.780 3395.220 111.180 3395.720 ;
        RECT 116.230 3395.220 116.630 3395.720 ;
        RECT 121.680 3395.220 122.080 3395.720 ;
        RECT 131.280 3395.220 131.680 3395.720 ;
        RECT 140.780 3395.220 141.180 3395.720 ;
        RECT 146.230 3395.220 146.630 3395.720 ;
        RECT 151.680 3395.220 152.080 3395.720 ;
        RECT 76.030 3394.070 76.430 3394.570 ;
        RECT 90.980 3394.070 91.380 3394.570 ;
        RECT 106.030 3394.070 106.430 3394.570 ;
        RECT 120.980 3394.070 121.380 3394.570 ;
        RECT 136.030 3394.070 136.430 3394.570 ;
        RECT 150.980 3394.070 151.380 3394.570 ;
        RECT 68.080 3393.570 75.080 3394.070 ;
        RECT 64.180 3349.370 65.180 3377.070 ;
        RECT 68.080 3366.720 68.580 3393.570 ;
        RECT 74.580 3390.470 75.080 3393.570 ;
        RECT 76.030 3393.570 105.080 3394.070 ;
        RECT 76.030 3393.170 76.430 3393.570 ;
        RECT 83.380 3390.470 83.880 3393.570 ;
        RECT 90.980 3393.170 91.380 3393.570 ;
        RECT 85.530 3392.520 85.930 3392.870 ;
        RECT 96.430 3392.520 96.830 3392.870 ;
        RECT 85.530 3392.020 96.830 3392.520 ;
        RECT 85.530 3391.670 85.930 3392.020 ;
        RECT 88.230 3390.470 88.730 3392.020 ;
        RECT 96.430 3391.670 96.830 3392.020 ;
        RECT 104.580 3390.470 105.080 3393.570 ;
        RECT 106.030 3393.570 135.080 3394.070 ;
        RECT 106.030 3393.170 106.430 3393.570 ;
        RECT 113.380 3390.470 113.880 3393.570 ;
        RECT 120.980 3393.170 121.380 3393.570 ;
        RECT 115.530 3392.520 115.930 3392.870 ;
        RECT 126.430 3392.520 126.830 3392.870 ;
        RECT 115.530 3392.020 126.830 3392.520 ;
        RECT 115.530 3391.670 115.930 3392.020 ;
        RECT 118.230 3390.470 118.730 3392.020 ;
        RECT 126.430 3391.670 126.830 3392.020 ;
        RECT 134.580 3390.470 135.080 3393.570 ;
        RECT 136.030 3393.570 165.980 3394.070 ;
        RECT 136.030 3393.170 136.430 3393.570 ;
        RECT 143.380 3390.470 143.880 3393.570 ;
        RECT 150.980 3393.170 151.380 3393.570 ;
        RECT 145.530 3392.520 145.930 3392.870 ;
        RECT 156.430 3392.520 156.830 3392.870 ;
        RECT 145.530 3392.020 156.830 3392.520 ;
        RECT 145.530 3391.670 145.930 3392.020 ;
        RECT 148.230 3390.470 148.730 3392.020 ;
        RECT 156.430 3391.670 156.830 3392.020 ;
        RECT 73.180 3389.820 78.080 3390.470 ;
        RECT 83.030 3389.820 84.230 3390.470 ;
        RECT 87.880 3389.820 89.080 3390.470 ;
        RECT 93.580 3390.370 98.480 3390.470 ;
        RECT 92.730 3389.870 98.480 3390.370 ;
        RECT 92.730 3387.720 93.230 3389.870 ;
        RECT 93.580 3389.820 98.480 3389.870 ;
        RECT 103.180 3389.820 108.080 3390.470 ;
        RECT 113.030 3389.820 114.230 3390.470 ;
        RECT 117.880 3389.820 119.080 3390.470 ;
        RECT 123.580 3390.370 128.480 3390.470 ;
        RECT 122.730 3389.870 128.480 3390.370 ;
        RECT 69.580 3387.220 93.230 3387.720 ;
        RECT 96.430 3387.720 96.830 3388.020 ;
        RECT 122.730 3387.720 123.230 3389.870 ;
        RECT 123.580 3389.820 128.480 3389.870 ;
        RECT 133.180 3389.820 138.080 3390.470 ;
        RECT 143.030 3389.820 144.230 3390.470 ;
        RECT 147.880 3389.820 149.080 3390.470 ;
        RECT 153.580 3390.370 158.480 3390.470 ;
        RECT 152.730 3389.870 158.480 3390.370 ;
        RECT 96.430 3387.220 123.230 3387.720 ;
        RECT 126.430 3387.720 126.830 3388.020 ;
        RECT 152.730 3387.720 153.230 3389.870 ;
        RECT 153.580 3389.820 158.480 3389.870 ;
        RECT 126.430 3387.220 153.230 3387.720 ;
        RECT 156.430 3387.720 156.830 3388.020 ;
        RECT 156.430 3387.220 163.080 3387.720 ;
        RECT 69.580 3373.070 70.080 3387.220 ;
        RECT 96.430 3386.820 96.830 3387.220 ;
        RECT 126.430 3386.820 126.830 3387.220 ;
        RECT 156.430 3386.820 156.830 3387.220 ;
        RECT 71.280 3383.320 71.680 3386.070 ;
        RECT 80.780 3383.320 81.180 3386.070 ;
        RECT 86.230 3383.320 86.630 3386.070 ;
        RECT 91.680 3383.320 92.080 3386.070 ;
        RECT 101.280 3383.320 101.680 3386.070 ;
        RECT 110.780 3383.320 111.180 3386.070 ;
        RECT 116.230 3383.320 116.630 3386.070 ;
        RECT 121.680 3383.320 122.080 3386.070 ;
        RECT 131.280 3383.320 131.680 3386.070 ;
        RECT 140.780 3383.320 141.180 3386.070 ;
        RECT 146.230 3383.320 146.630 3386.070 ;
        RECT 151.680 3383.320 152.080 3386.070 ;
        RECT 71.280 3382.820 152.080 3383.320 ;
        RECT 93.630 3378.670 97.830 3379.170 ;
        RECT 93.730 3377.970 94.230 3378.670 ;
        RECT 93.720 3377.490 96.020 3377.970 ;
        RECT 72.030 3376.070 93.430 3377.070 ;
        RECT 96.280 3376.870 96.680 3378.670 ;
        RECT 95.530 3376.470 96.130 3376.770 ;
        RECT 97.330 3376.470 97.830 3378.670 ;
        RECT 95.530 3376.170 97.830 3376.470 ;
        RECT 95.480 3375.820 95.930 3375.920 ;
        RECT 92.530 3375.520 95.930 3375.820 ;
        RECT 92.530 3373.070 93.030 3375.520 ;
        RECT 95.480 3375.470 95.930 3375.520 ;
        RECT 96.280 3375.720 96.680 3375.870 ;
        RECT 99.230 3375.720 99.730 3382.820 ;
        RECT 103.150 3380.870 105.255 3381.250 ;
        RECT 110.080 3379.770 110.580 3382.820 ;
        RECT 109.230 3379.700 110.580 3379.770 ;
        RECT 103.150 3379.320 105.255 3379.700 ;
        RECT 107.305 3379.320 110.580 3379.700 ;
        RECT 109.230 3379.220 110.580 3379.320 ;
        RECT 96.280 3375.420 99.730 3375.720 ;
        RECT 96.280 3375.370 96.680 3375.420 ;
        RECT 93.720 3375.070 96.020 3375.250 ;
        RECT 99.230 3375.070 99.730 3375.420 ;
        RECT 93.720 3374.770 99.730 3375.070 ;
        RECT 110.080 3377.470 110.580 3379.220 ;
        RECT 151.580 3377.470 152.080 3382.820 ;
        RECT 110.080 3376.970 160.880 3377.470 ;
        RECT 110.080 3374.220 110.480 3376.970 ;
        RECT 115.530 3374.220 115.930 3376.970 ;
        RECT 120.980 3374.220 121.380 3376.970 ;
        RECT 130.480 3374.220 130.880 3376.970 ;
        RECT 140.080 3374.220 140.480 3376.970 ;
        RECT 145.530 3374.220 145.930 3376.970 ;
        RECT 150.980 3374.220 151.380 3376.970 ;
        RECT 160.480 3374.220 160.880 3376.970 ;
        RECT 105.330 3373.070 105.730 3373.470 ;
        RECT 135.330 3373.070 135.730 3373.470 ;
        RECT 162.080 3373.070 163.080 3387.220 ;
        RECT 69.580 3372.570 105.730 3373.070 ;
        RECT 105.330 3372.270 105.730 3372.570 ;
        RECT 108.930 3372.570 135.730 3373.070 ;
        RECT 103.680 3370.420 108.580 3370.470 ;
        RECT 108.930 3370.420 109.430 3372.570 ;
        RECT 135.330 3372.270 135.730 3372.570 ;
        RECT 138.930 3372.570 163.080 3373.070 ;
        RECT 103.680 3369.920 109.430 3370.420 ;
        RECT 103.680 3369.820 108.580 3369.920 ;
        RECT 113.080 3369.820 114.280 3370.470 ;
        RECT 117.930 3369.820 119.130 3370.470 ;
        RECT 124.080 3369.820 128.980 3370.470 ;
        RECT 133.680 3370.420 138.580 3370.470 ;
        RECT 138.930 3370.420 139.430 3372.570 ;
        RECT 133.680 3369.920 139.430 3370.420 ;
        RECT 133.680 3369.820 138.580 3369.920 ;
        RECT 143.080 3369.820 144.280 3370.470 ;
        RECT 147.930 3369.820 149.130 3370.470 ;
        RECT 154.080 3369.820 158.980 3370.470 ;
        RECT 105.330 3368.270 105.730 3368.620 ;
        RECT 113.430 3368.270 113.930 3369.820 ;
        RECT 116.230 3368.270 116.630 3368.620 ;
        RECT 105.330 3367.770 116.630 3368.270 ;
        RECT 105.330 3367.420 105.730 3367.770 ;
        RECT 116.230 3367.420 116.630 3367.770 ;
        RECT 110.780 3366.720 111.180 3367.120 ;
        RECT 118.280 3366.720 118.780 3369.820 ;
        RECT 125.730 3366.720 126.130 3367.120 ;
        RECT 68.080 3366.220 126.130 3366.720 ;
        RECT 127.080 3366.720 127.580 3369.820 ;
        RECT 135.330 3368.270 135.730 3368.620 ;
        RECT 143.430 3368.270 143.930 3369.820 ;
        RECT 146.230 3368.270 146.630 3368.620 ;
        RECT 135.330 3367.770 146.630 3368.270 ;
        RECT 135.330 3367.420 135.730 3367.770 ;
        RECT 146.230 3367.420 146.630 3367.770 ;
        RECT 140.780 3366.720 141.180 3367.120 ;
        RECT 148.280 3366.720 148.780 3369.820 ;
        RECT 155.730 3366.720 156.130 3367.120 ;
        RECT 127.080 3366.220 156.130 3366.720 ;
        RECT 157.080 3366.720 157.580 3369.820 ;
        RECT 164.980 3366.720 165.980 3393.570 ;
        RECT 157.080 3366.220 165.980 3366.720 ;
        RECT 68.080 3354.570 68.580 3366.220 ;
        RECT 110.780 3365.720 111.180 3366.220 ;
        RECT 125.730 3365.720 126.130 3366.220 ;
        RECT 140.780 3365.720 141.180 3366.220 ;
        RECT 155.730 3365.720 156.130 3366.220 ;
        RECT 110.080 3364.570 110.480 3365.070 ;
        RECT 115.530 3364.570 115.930 3365.070 ;
        RECT 120.980 3364.570 121.380 3365.070 ;
        RECT 130.480 3364.570 130.880 3365.070 ;
        RECT 140.080 3364.570 140.480 3365.070 ;
        RECT 145.530 3364.570 145.930 3365.070 ;
        RECT 150.980 3364.570 151.380 3365.070 ;
        RECT 160.480 3364.570 160.880 3365.070 ;
        RECT 70.780 3356.140 72.780 3362.170 ;
        RECT 76.580 3356.140 78.580 3362.170 ;
        RECT 82.630 3356.140 84.630 3362.170 ;
        RECT 87.630 3361.770 88.180 3364.570 ;
        RECT 87.630 3361.170 108.680 3361.770 ;
        RECT 68.970 3355.660 85.720 3356.140 ;
        RECT 70.780 3355.640 72.480 3355.660 ;
        RECT 82.030 3355.640 83.880 3355.660 ;
        RECT 87.380 3355.640 88.180 3355.990 ;
        RECT 71.430 3355.040 71.830 3355.640 ;
        RECT 72.960 3355.120 73.250 3355.165 ;
        RECT 74.820 3355.120 75.110 3355.165 ;
        RECT 77.600 3355.120 77.890 3355.165 ;
        RECT 72.960 3354.980 77.890 3355.120 ;
        RECT 72.960 3354.935 73.250 3354.980 ;
        RECT 74.820 3354.935 75.110 3354.980 ;
        RECT 77.600 3354.935 77.890 3354.980 ;
        RECT 84.930 3354.940 87.230 3355.290 ;
        RECT 68.080 3354.170 68.880 3354.570 ;
        RECT 71.430 3354.290 74.580 3354.690 ;
        RECT 77.600 3354.440 77.890 3354.485 ;
        RECT 75.355 3354.300 77.890 3354.440 ;
        RECT 68.380 3353.440 68.780 3353.940 ;
        RECT 68.380 3353.420 69.080 3353.440 ;
        RECT 68.380 3352.940 70.810 3353.420 ;
        RECT 68.430 3350.930 69.180 3350.940 ;
        RECT 68.430 3350.450 70.500 3350.930 ;
        RECT 68.430 3350.440 69.180 3350.450 ;
        RECT 68.430 3349.990 68.830 3350.440 ;
        RECT 64.180 3348.970 69.580 3349.370 ;
        RECT 70.130 3349.340 70.580 3349.390 ;
        RECT 69.730 3348.990 70.580 3349.340 ;
        RECT 64.180 3317.720 65.180 3348.970 ;
        RECT 70.130 3348.940 70.580 3348.990 ;
        RECT 68.430 3348.240 68.830 3348.740 ;
        RECT 68.430 3348.210 69.130 3348.240 ;
        RECT 68.430 3347.730 70.500 3348.210 ;
        RECT 68.430 3347.690 69.130 3347.730 ;
        RECT 71.430 3347.440 71.780 3354.290 ;
        RECT 75.355 3354.145 75.570 3354.300 ;
        RECT 77.600 3354.255 77.890 3354.300 ;
        RECT 73.420 3354.100 73.710 3354.145 ;
        RECT 75.280 3354.100 75.570 3354.145 ;
        RECT 76.200 3354.140 76.490 3354.145 ;
        RECT 73.420 3353.960 75.570 3354.100 ;
        RECT 73.420 3353.915 73.710 3353.960 ;
        RECT 75.280 3353.915 75.570 3353.960 ;
        RECT 76.130 3354.100 76.630 3354.140 ;
        RECT 79.460 3354.100 79.750 3354.145 ;
        RECT 76.130 3353.960 79.750 3354.100 ;
        RECT 76.130 3353.690 76.630 3353.960 ;
        RECT 79.460 3353.915 79.750 3353.960 ;
        RECT 72.410 3352.940 82.070 3353.420 ;
        RECT 74.680 3347.890 75.030 3352.940 ;
        RECT 82.880 3351.690 83.230 3354.540 ;
        RECT 83.880 3352.940 85.720 3353.420 ;
        RECT 75.530 3351.340 83.230 3351.690 ;
        RECT 75.530 3349.690 75.880 3351.340 ;
        RECT 80.330 3350.460 81.730 3350.490 ;
        RECT 77.130 3349.990 83.550 3350.460 ;
        RECT 77.130 3349.980 80.350 3349.990 ;
        RECT 75.530 3349.340 78.430 3349.690 ;
        RECT 77.480 3348.490 77.830 3348.840 ;
        RECT 78.080 3348.790 78.430 3349.340 ;
        RECT 80.880 3349.240 81.280 3349.990 ;
        RECT 81.710 3349.980 83.550 3349.990 ;
        RECT 82.730 3348.920 83.030 3349.590 ;
        RECT 77.980 3348.540 78.530 3348.790 ;
        RECT 82.730 3348.530 84.630 3348.920 ;
        RECT 83.030 3348.520 84.630 3348.530 ;
        RECT 75.530 3348.140 77.830 3348.490 ;
        RECT 68.780 3347.140 71.780 3347.440 ;
        RECT 68.780 3344.990 69.130 3347.140 ;
        RECT 75.530 3346.440 75.880 3348.140 ;
        RECT 80.780 3347.740 81.280 3348.140 ;
        RECT 77.130 3347.260 83.550 3347.740 ;
        RECT 80.330 3347.240 81.730 3347.260 ;
        RECT 86.880 3346.640 87.230 3354.940 ;
        RECT 71.780 3346.090 75.880 3346.440 ;
        RECT 82.530 3346.290 87.230 3346.640 ;
        RECT 69.980 3345.290 71.360 3345.770 ;
        RECT 71.780 3345.040 72.130 3346.090 ;
        RECT 72.450 3345.290 82.110 3345.770 ;
        RECT 68.780 3344.640 70.830 3344.990 ;
        RECT 71.780 3344.640 73.230 3345.040 ;
        RECT 74.770 3344.750 75.060 3344.795 ;
        RECT 78.030 3344.750 78.530 3345.090 ;
        RECT 74.770 3344.610 78.530 3344.750 ;
        RECT 74.770 3344.565 75.060 3344.610 ;
        RECT 78.030 3344.590 78.530 3344.610 ;
        RECT 78.950 3344.750 79.240 3344.795 ;
        RECT 80.810 3344.750 81.100 3344.795 ;
        RECT 78.950 3344.610 81.100 3344.750 ;
        RECT 78.030 3344.565 78.320 3344.590 ;
        RECT 78.950 3344.565 79.240 3344.610 ;
        RECT 80.810 3344.565 81.100 3344.610 ;
        RECT 76.630 3344.410 76.920 3344.455 ;
        RECT 78.950 3344.410 79.165 3344.565 ;
        RECT 76.630 3344.270 79.165 3344.410 ;
        RECT 76.630 3344.225 76.920 3344.270 ;
        RECT 79.930 3344.240 80.330 3344.440 ;
        RECT 82.530 3344.240 82.880 3346.290 ;
        RECT 84.040 3345.290 85.880 3345.770 ;
        RECT 83.180 3344.890 83.680 3345.290 ;
        RECT 79.930 3343.940 82.880 3344.240 ;
        RECT 83.230 3344.190 84.880 3344.540 ;
        RECT 79.930 3343.890 81.130 3343.940 ;
        RECT 81.730 3343.890 82.880 3343.940 ;
        RECT 69.980 3343.040 71.360 3343.050 ;
        RECT 71.830 3343.040 72.230 3343.790 ;
        RECT 76.630 3343.730 76.920 3343.775 ;
        RECT 79.410 3343.730 79.700 3343.775 ;
        RECT 81.270 3343.730 81.560 3343.775 ;
        RECT 76.630 3343.590 81.560 3343.730 ;
        RECT 76.630 3343.545 76.920 3343.590 ;
        RECT 79.410 3343.545 79.700 3343.590 ;
        RECT 81.270 3343.545 81.560 3343.590 ;
        RECT 84.530 3343.390 84.880 3344.190 ;
        RECT 72.450 3343.040 82.110 3343.050 ;
        RECT 84.040 3343.040 85.880 3343.050 ;
        RECT 69.980 3342.590 85.880 3343.040 ;
        RECT 87.830 3342.940 88.180 3355.640 ;
        RECT 108.080 3350.470 108.680 3361.170 ;
        RECT 157.980 3360.170 164.980 3360.570 ;
        RECT 112.780 3358.820 113.180 3359.320 ;
        RECT 117.480 3358.720 117.880 3359.220 ;
        RECT 120.580 3358.720 120.980 3359.220 ;
        RECT 123.680 3358.820 124.080 3359.320 ;
        RECT 128.380 3358.820 128.780 3359.320 ;
        RECT 133.080 3358.720 133.480 3359.220 ;
        RECT 136.180 3358.720 136.580 3359.220 ;
        RECT 139.280 3358.820 139.680 3359.320 ;
        RECT 143.980 3358.820 144.380 3359.320 ;
        RECT 148.680 3358.720 149.080 3359.220 ;
        RECT 151.780 3358.720 152.180 3359.220 ;
        RECT 154.880 3358.820 155.280 3359.320 ;
        RECT 115.080 3358.270 115.480 3358.470 ;
        RECT 122.880 3358.270 123.280 3358.470 ;
        RECT 115.080 3358.070 123.280 3358.270 ;
        RECT 130.680 3358.270 131.080 3358.470 ;
        RECT 138.480 3358.270 138.880 3358.470 ;
        RECT 130.680 3358.070 138.880 3358.270 ;
        RECT 146.280 3358.270 146.680 3358.470 ;
        RECT 154.080 3358.270 154.480 3358.470 ;
        RECT 146.280 3358.070 154.480 3358.270 ;
        RECT 110.080 3357.670 114.530 3358.070 ;
        RECT 115.080 3357.870 130.130 3358.070 ;
        RECT 115.080 3357.670 115.480 3357.870 ;
        RECT 108.080 3349.970 109.030 3350.470 ;
        RECT 107.930 3348.520 108.730 3348.920 ;
        RECT 90.180 3345.470 91.880 3345.970 ;
        RECT 87.430 3342.590 88.180 3342.940 ;
        RECT 69.980 3342.570 71.360 3342.590 ;
        RECT 72.450 3342.570 82.110 3342.590 ;
        RECT 84.040 3342.570 85.880 3342.590 ;
        RECT 89.980 3339.220 91.980 3345.470 ;
        RECT 97.580 3344.120 98.780 3344.720 ;
        RECT 98.180 3342.970 98.780 3344.120 ;
        RECT 66.580 3336.640 95.250 3337.120 ;
        RECT 66.580 3336.620 70.880 3336.640 ;
        RECT 74.430 3336.620 74.930 3336.640 ;
        RECT 78.530 3336.620 79.030 3336.640 ;
        RECT 82.630 3336.620 83.380 3336.640 ;
        RECT 87.030 3336.620 87.480 3336.640 ;
        RECT 91.130 3336.620 91.580 3336.640 ;
        RECT 66.580 3333.120 68.580 3336.620 ;
        RECT 82.880 3335.970 83.280 3336.620 ;
        RECT 70.860 3335.670 71.560 3335.790 ;
        RECT 69.330 3335.320 71.560 3335.670 ;
        RECT 69.330 3333.670 70.330 3335.320 ;
        RECT 70.860 3335.220 71.560 3335.320 ;
        RECT 82.830 3334.420 83.140 3334.910 ;
        RECT 74.430 3334.400 74.880 3334.420 ;
        RECT 78.530 3334.400 78.980 3334.420 ;
        RECT 82.630 3334.400 83.380 3334.420 ;
        RECT 87.030 3334.400 87.480 3334.420 ;
        RECT 91.130 3334.400 91.580 3334.420 ;
        RECT 70.770 3333.920 95.250 3334.400 ;
        RECT 69.330 3333.320 74.180 3333.670 ;
        RECT 66.580 3332.640 72.610 3333.120 ;
        RECT 66.580 3332.620 70.880 3332.640 ;
        RECT 71.800 3331.610 72.100 3332.460 ;
        RECT 73.030 3331.970 73.430 3332.470 ;
        RECT 70.830 3331.520 71.230 3331.570 ;
        RECT 69.230 3331.170 71.230 3331.520 ;
        RECT 71.810 3331.510 72.100 3331.610 ;
        RECT 73.830 3331.820 74.180 3333.320 ;
        RECT 74.570 3332.640 87.850 3333.120 ;
        RECT 81.930 3332.620 83.830 3332.640 ;
        RECT 85.180 3332.620 86.480 3332.640 ;
        RECT 86.980 3332.220 87.380 3332.370 ;
        RECT 88.480 3332.220 90.280 3332.320 ;
        RECT 75.140 3332.100 75.430 3332.145 ;
        RECT 77.240 3332.100 77.530 3332.145 ;
        RECT 78.810 3332.100 79.100 3332.145 ;
        RECT 75.140 3331.960 79.100 3332.100 ;
        RECT 75.140 3331.915 75.430 3331.960 ;
        RECT 77.240 3331.915 77.530 3331.960 ;
        RECT 78.810 3331.915 79.100 3331.960 ;
        RECT 86.980 3331.870 90.280 3332.220 ;
        RECT 73.830 3331.780 74.980 3331.820 ;
        RECT 71.810 3331.210 73.690 3331.510 ;
        RECT 73.830 3331.470 74.990 3331.780 ;
        RECT 75.535 3331.760 75.825 3331.805 ;
        RECT 76.725 3331.760 77.015 3331.805 ;
        RECT 79.245 3331.760 79.535 3331.805 ;
        RECT 75.535 3331.620 79.535 3331.760 ;
        RECT 88.480 3331.720 90.280 3331.870 ;
        RECT 75.535 3331.575 75.825 3331.620 ;
        RECT 76.725 3331.575 77.015 3331.620 ;
        RECT 79.245 3331.575 79.535 3331.620 ;
        RECT 69.230 3326.270 69.630 3331.170 ;
        RECT 70.830 3331.120 71.230 3331.170 ;
        RECT 72.780 3330.420 73.180 3331.020 ;
        RECT 73.460 3330.920 73.690 3331.210 ;
        RECT 74.640 3331.130 74.990 3331.470 ;
        RECT 75.920 3330.920 76.200 3331.210 ;
        RECT 86.180 3331.170 86.930 3331.520 ;
        RECT 86.180 3331.070 86.480 3331.170 ;
        RECT 73.460 3330.620 76.200 3330.920 ;
        RECT 84.430 3330.770 86.480 3331.070 ;
        RECT 90.590 3330.420 91.065 3333.920 ;
        RECT 98.185 3332.920 98.780 3342.970 ;
        RECT 98.180 3332.320 98.780 3332.920 ;
        RECT 97.580 3331.720 98.780 3332.320 ;
        RECT 108.330 3332.470 108.730 3348.520 ;
        RECT 110.080 3342.470 110.580 3357.670 ;
        RECT 114.130 3355.920 114.530 3357.670 ;
        RECT 117.480 3355.970 117.880 3357.870 ;
        RECT 122.880 3357.670 130.130 3357.870 ;
        RECT 130.680 3357.870 145.730 3358.070 ;
        RECT 130.680 3357.670 131.080 3357.870 ;
        RECT 125.980 3357.070 126.380 3357.270 ;
        RECT 122.030 3356.620 126.380 3357.070 ;
        RECT 122.030 3355.970 122.480 3356.620 ;
        RECT 125.980 3356.470 126.380 3356.620 ;
        RECT 114.130 3355.470 116.180 3355.920 ;
        RECT 117.480 3355.470 119.780 3355.970 ;
        RECT 121.680 3355.470 122.630 3355.970 ;
        RECT 129.730 3355.920 130.130 3357.670 ;
        RECT 133.080 3355.970 133.480 3357.870 ;
        RECT 138.480 3357.670 145.730 3357.870 ;
        RECT 146.280 3357.870 163.480 3358.070 ;
        RECT 146.280 3357.670 146.680 3357.870 ;
        RECT 141.580 3357.070 141.980 3357.270 ;
        RECT 137.630 3356.620 141.980 3357.070 ;
        RECT 137.630 3355.970 138.080 3356.620 ;
        RECT 141.580 3356.470 141.980 3356.620 ;
        RECT 123.680 3355.470 127.080 3355.920 ;
        RECT 129.730 3355.470 131.780 3355.920 ;
        RECT 133.080 3355.470 135.380 3355.970 ;
        RECT 137.280 3355.470 138.230 3355.970 ;
        RECT 145.330 3355.920 145.730 3357.670 ;
        RECT 148.680 3355.970 149.080 3357.870 ;
        RECT 154.080 3357.670 163.480 3357.870 ;
        RECT 157.180 3357.070 157.580 3357.270 ;
        RECT 153.230 3356.620 157.580 3357.070 ;
        RECT 153.230 3355.970 153.680 3356.620 ;
        RECT 157.180 3356.470 157.580 3356.620 ;
        RECT 139.280 3355.470 142.680 3355.920 ;
        RECT 145.330 3355.470 147.380 3355.920 ;
        RECT 148.680 3355.470 150.980 3355.970 ;
        RECT 152.880 3355.470 153.830 3355.970 ;
        RECT 154.880 3355.470 158.280 3355.920 ;
        RECT 123.680 3354.370 124.080 3355.470 ;
        RECT 111.580 3353.970 124.080 3354.370 ;
        RECT 125.980 3354.370 126.380 3354.770 ;
        RECT 139.280 3354.370 139.680 3355.470 ;
        RECT 125.980 3353.970 139.680 3354.370 ;
        RECT 141.580 3354.370 141.980 3354.770 ;
        RECT 154.880 3354.370 155.280 3355.470 ;
        RECT 141.580 3353.970 155.280 3354.370 ;
        RECT 157.180 3354.370 157.580 3354.770 ;
        RECT 157.180 3353.970 161.980 3354.370 ;
        RECT 111.580 3346.170 112.080 3353.970 ;
        RECT 112.780 3353.120 113.180 3353.620 ;
        RECT 117.480 3353.120 117.880 3353.620 ;
        RECT 120.580 3353.120 120.980 3353.620 ;
        RECT 123.680 3353.120 124.080 3353.620 ;
        RECT 125.980 3353.570 126.380 3353.970 ;
        RECT 128.380 3353.120 128.780 3353.620 ;
        RECT 133.080 3353.120 133.480 3353.620 ;
        RECT 136.180 3353.120 136.580 3353.620 ;
        RECT 139.280 3353.120 139.680 3353.620 ;
        RECT 141.580 3353.570 141.980 3353.970 ;
        RECT 143.980 3353.120 144.380 3353.620 ;
        RECT 148.680 3353.120 149.080 3353.620 ;
        RECT 151.780 3353.120 152.180 3353.620 ;
        RECT 154.880 3353.120 155.280 3353.620 ;
        RECT 157.180 3353.570 157.580 3353.970 ;
        RECT 115.280 3349.370 123.780 3349.820 ;
        RECT 119.980 3348.650 120.280 3349.370 ;
        RECT 120.620 3349.340 122.920 3349.370 ;
        RECT 113.580 3347.820 121.180 3348.370 ;
        RECT 123.430 3348.170 123.780 3349.370 ;
        RECT 127.230 3348.270 127.630 3348.820 ;
        RECT 122.580 3347.820 123.780 3348.170 ;
        RECT 125.780 3347.870 128.180 3348.270 ;
        RECT 120.070 3347.070 120.380 3347.550 ;
        RECT 120.620 3347.070 122.920 3347.100 ;
        RECT 125.780 3347.070 126.280 3347.870 ;
        RECT 120.030 3346.620 126.280 3347.070 ;
        RECT 128.830 3346.170 129.230 3346.570 ;
        RECT 131.130 3346.520 131.530 3347.020 ;
        RECT 134.230 3346.520 134.630 3347.020 ;
        RECT 137.330 3346.520 137.730 3347.020 ;
        RECT 142.030 3346.520 142.430 3347.020 ;
        RECT 144.430 3346.170 144.830 3346.570 ;
        RECT 146.730 3346.520 147.130 3347.020 ;
        RECT 149.830 3346.520 150.230 3347.020 ;
        RECT 152.930 3346.520 153.330 3347.020 ;
        RECT 157.630 3346.520 158.030 3347.020 ;
        RECT 161.480 3346.170 161.980 3353.970 ;
        RECT 111.580 3345.770 129.230 3346.170 ;
        RECT 128.830 3345.370 129.230 3345.770 ;
        RECT 131.130 3345.770 144.830 3346.170 ;
        RECT 131.130 3344.670 131.530 3345.770 ;
        RECT 144.430 3345.370 144.830 3345.770 ;
        RECT 146.730 3345.770 161.980 3346.170 ;
        RECT 146.730 3344.670 147.130 3345.770 ;
        RECT 128.130 3344.220 131.530 3344.670 ;
        RECT 132.580 3344.170 133.530 3344.670 ;
        RECT 135.430 3344.170 137.730 3344.670 ;
        RECT 139.030 3344.220 141.080 3344.670 ;
        RECT 143.730 3344.220 147.130 3344.670 ;
        RECT 128.830 3343.520 129.230 3343.670 ;
        RECT 132.730 3343.520 133.180 3344.170 ;
        RECT 128.830 3343.070 133.180 3343.520 ;
        RECT 128.830 3342.870 129.230 3343.070 ;
        RECT 110.080 3342.270 132.330 3342.470 ;
        RECT 137.330 3342.270 137.730 3344.170 ;
        RECT 140.680 3342.470 141.080 3344.220 ;
        RECT 148.180 3344.170 149.130 3344.670 ;
        RECT 151.030 3344.170 153.330 3344.670 ;
        RECT 154.630 3344.220 156.680 3344.670 ;
        RECT 144.430 3343.520 144.830 3343.670 ;
        RECT 148.330 3343.520 148.780 3344.170 ;
        RECT 144.430 3343.070 148.780 3343.520 ;
        RECT 144.430 3342.870 144.830 3343.070 ;
        RECT 139.730 3342.270 140.130 3342.470 ;
        RECT 110.080 3342.070 140.130 3342.270 ;
        RECT 140.680 3342.270 147.930 3342.470 ;
        RECT 152.930 3342.270 153.330 3344.170 ;
        RECT 156.280 3342.470 156.680 3344.220 ;
        RECT 162.980 3342.470 163.480 3357.670 ;
        RECT 155.330 3342.270 155.730 3342.470 ;
        RECT 140.680 3342.070 155.730 3342.270 ;
        RECT 156.280 3342.070 163.480 3342.470 ;
        RECT 125.280 3336.270 125.680 3342.070 ;
        RECT 131.930 3341.870 140.130 3342.070 ;
        RECT 131.930 3341.670 132.330 3341.870 ;
        RECT 139.730 3341.670 140.130 3341.870 ;
        RECT 147.530 3341.870 155.730 3342.070 ;
        RECT 147.530 3341.670 147.930 3341.870 ;
        RECT 155.330 3341.670 155.730 3341.870 ;
        RECT 131.130 3340.820 131.530 3341.320 ;
        RECT 134.230 3340.920 134.630 3341.420 ;
        RECT 137.330 3340.920 137.730 3341.420 ;
        RECT 142.030 3340.820 142.430 3341.320 ;
        RECT 146.730 3340.820 147.130 3341.320 ;
        RECT 149.830 3340.920 150.230 3341.420 ;
        RECT 152.930 3340.920 153.330 3341.420 ;
        RECT 157.630 3340.820 158.030 3341.320 ;
        RECT 164.480 3339.970 164.980 3360.170 ;
        RECT 170.130 3347.870 171.230 3348.370 ;
        RECT 156.830 3339.570 164.980 3339.970 ;
        RECT 143.980 3337.620 144.430 3338.920 ;
        RECT 143.380 3337.170 144.430 3337.620 ;
        RECT 125.280 3335.870 136.630 3336.270 ;
        RECT 138.220 3335.940 140.060 3336.420 ;
        RECT 136.230 3334.820 136.630 3335.870 ;
        RECT 136.230 3334.810 138.330 3334.820 ;
        RECT 136.230 3334.450 138.660 3334.810 ;
        RECT 139.280 3334.770 139.530 3335.770 ;
        RECT 140.330 3335.020 140.630 3335.520 ;
        RECT 140.930 3334.770 145.530 3334.920 ;
        RECT 139.280 3334.570 145.530 3334.770 ;
        RECT 139.365 3334.560 145.530 3334.570 ;
        RECT 136.230 3334.420 138.330 3334.450 ;
        RECT 140.930 3334.420 145.530 3334.560 ;
        RECT 138.220 3333.670 140.060 3333.700 ;
        RECT 140.330 3333.670 140.630 3334.270 ;
        RECT 137.830 3333.220 140.630 3333.670 ;
        RECT 108.330 3332.070 110.780 3332.470 ;
        RECT 98.180 3331.120 98.780 3331.720 ;
        RECT 72.580 3330.400 74.580 3330.420 ;
        RECT 81.930 3330.400 83.830 3330.420 ;
        RECT 85.180 3330.400 86.480 3330.420 ;
        RECT 87.780 3330.400 91.065 3330.420 ;
        RECT 70.770 3329.920 91.065 3330.400 ;
        RECT 70.780 3328.720 72.780 3329.920 ;
        RECT 79.430 3328.720 81.430 3329.920 ;
        RECT 88.630 3328.720 90.630 3329.920 ;
        RECT 69.230 3325.870 90.030 3326.270 ;
        RECT 68.970 3324.010 85.720 3324.490 ;
        RECT 70.780 3323.990 72.480 3324.010 ;
        RECT 82.030 3323.990 83.880 3324.010 ;
        RECT 87.380 3323.990 88.180 3324.340 ;
        RECT 71.430 3323.390 71.830 3323.990 ;
        RECT 72.960 3323.470 73.250 3323.515 ;
        RECT 74.820 3323.470 75.110 3323.515 ;
        RECT 77.600 3323.470 77.890 3323.515 ;
        RECT 72.960 3323.330 77.890 3323.470 ;
        RECT 72.960 3323.285 73.250 3323.330 ;
        RECT 74.820 3323.285 75.110 3323.330 ;
        RECT 77.600 3323.285 77.890 3323.330 ;
        RECT 84.930 3323.290 87.230 3323.640 ;
        RECT 66.980 3322.520 67.780 3322.920 ;
        RECT 71.430 3322.640 74.580 3323.040 ;
        RECT 77.600 3322.790 77.890 3322.835 ;
        RECT 75.355 3322.650 77.890 3322.790 ;
        RECT 64.180 3317.320 65.380 3317.720 ;
        RECT 64.180 3315.420 65.180 3317.320 ;
        RECT 66.980 3306.520 67.380 3322.520 ;
        RECT 68.380 3321.790 68.780 3322.290 ;
        RECT 68.380 3321.770 69.080 3321.790 ;
        RECT 68.380 3321.290 70.810 3321.770 ;
        RECT 68.380 3320.770 70.780 3321.290 ;
        RECT 68.430 3319.280 69.180 3319.290 ;
        RECT 68.430 3318.800 70.500 3319.280 ;
        RECT 68.430 3318.790 69.180 3318.800 ;
        RECT 68.430 3318.340 68.830 3318.790 ;
        RECT 67.680 3317.320 69.580 3317.720 ;
        RECT 70.130 3317.690 70.580 3317.740 ;
        RECT 69.730 3317.340 70.580 3317.690 ;
        RECT 70.130 3317.290 70.580 3317.340 ;
        RECT 68.430 3316.590 68.830 3317.090 ;
        RECT 68.430 3316.560 69.130 3316.590 ;
        RECT 68.430 3316.080 70.500 3316.560 ;
        RECT 68.430 3316.040 69.130 3316.080 ;
        RECT 71.430 3315.790 71.780 3322.640 ;
        RECT 75.355 3322.495 75.570 3322.650 ;
        RECT 77.600 3322.605 77.890 3322.650 ;
        RECT 73.420 3322.450 73.710 3322.495 ;
        RECT 75.280 3322.450 75.570 3322.495 ;
        RECT 76.200 3322.490 76.490 3322.495 ;
        RECT 73.420 3322.310 75.570 3322.450 ;
        RECT 73.420 3322.265 73.710 3322.310 ;
        RECT 75.280 3322.265 75.570 3322.310 ;
        RECT 76.130 3322.450 76.630 3322.490 ;
        RECT 79.460 3322.450 79.750 3322.495 ;
        RECT 76.130 3322.310 79.750 3322.450 ;
        RECT 76.130 3322.040 76.630 3322.310 ;
        RECT 79.460 3322.265 79.750 3322.310 ;
        RECT 72.410 3321.290 82.070 3321.770 ;
        RECT 74.680 3316.240 75.030 3321.290 ;
        RECT 82.880 3320.040 83.230 3322.890 ;
        RECT 83.880 3321.290 85.720 3321.770 ;
        RECT 75.530 3319.690 83.230 3320.040 ;
        RECT 75.530 3318.040 75.880 3319.690 ;
        RECT 80.330 3318.810 81.730 3318.840 ;
        RECT 77.130 3318.340 83.550 3318.810 ;
        RECT 77.130 3318.330 80.350 3318.340 ;
        RECT 75.530 3317.690 78.430 3318.040 ;
        RECT 77.480 3316.840 77.830 3317.190 ;
        RECT 78.080 3317.140 78.430 3317.690 ;
        RECT 80.880 3317.590 81.280 3318.340 ;
        RECT 81.710 3318.330 83.550 3318.340 ;
        RECT 82.730 3317.270 83.030 3317.940 ;
        RECT 77.980 3316.890 78.530 3317.140 ;
        RECT 82.730 3316.880 85.680 3317.270 ;
        RECT 83.030 3316.870 85.680 3316.880 ;
        RECT 75.530 3316.490 77.830 3316.840 ;
        RECT 68.780 3315.490 71.780 3315.790 ;
        RECT 68.780 3313.340 69.130 3315.490 ;
        RECT 75.530 3314.790 75.880 3316.490 ;
        RECT 80.780 3316.090 81.280 3316.490 ;
        RECT 77.130 3315.610 83.550 3316.090 ;
        RECT 80.330 3315.590 81.730 3315.610 ;
        RECT 86.880 3314.990 87.230 3323.290 ;
        RECT 71.780 3314.440 75.880 3314.790 ;
        RECT 82.530 3314.640 87.230 3314.990 ;
        RECT 69.980 3313.640 71.360 3314.120 ;
        RECT 71.780 3313.390 72.130 3314.440 ;
        RECT 72.450 3313.640 82.110 3314.120 ;
        RECT 68.780 3312.990 70.830 3313.340 ;
        RECT 71.780 3312.990 73.230 3313.390 ;
        RECT 74.770 3313.100 75.060 3313.145 ;
        RECT 78.030 3313.100 78.530 3313.440 ;
        RECT 74.770 3312.960 78.530 3313.100 ;
        RECT 74.770 3312.915 75.060 3312.960 ;
        RECT 78.030 3312.940 78.530 3312.960 ;
        RECT 78.950 3313.100 79.240 3313.145 ;
        RECT 80.810 3313.100 81.100 3313.145 ;
        RECT 78.950 3312.960 81.100 3313.100 ;
        RECT 78.030 3312.915 78.320 3312.940 ;
        RECT 78.950 3312.915 79.240 3312.960 ;
        RECT 80.810 3312.915 81.100 3312.960 ;
        RECT 76.630 3312.760 76.920 3312.805 ;
        RECT 78.950 3312.760 79.165 3312.915 ;
        RECT 76.630 3312.620 79.165 3312.760 ;
        RECT 76.630 3312.575 76.920 3312.620 ;
        RECT 79.930 3312.590 80.330 3312.790 ;
        RECT 82.530 3312.590 82.880 3314.640 ;
        RECT 84.040 3313.640 85.880 3314.120 ;
        RECT 83.180 3313.240 83.680 3313.640 ;
        RECT 79.930 3312.290 82.880 3312.590 ;
        RECT 83.230 3312.540 84.880 3312.890 ;
        RECT 79.930 3312.240 81.130 3312.290 ;
        RECT 81.730 3312.240 82.880 3312.290 ;
        RECT 69.980 3311.390 71.360 3311.400 ;
        RECT 71.830 3311.390 72.230 3312.140 ;
        RECT 76.630 3312.080 76.920 3312.125 ;
        RECT 79.410 3312.080 79.700 3312.125 ;
        RECT 81.270 3312.080 81.560 3312.125 ;
        RECT 76.630 3311.940 81.560 3312.080 ;
        RECT 76.630 3311.895 76.920 3311.940 ;
        RECT 79.410 3311.895 79.700 3311.940 ;
        RECT 81.270 3311.895 81.560 3311.940 ;
        RECT 84.530 3311.740 84.880 3312.540 ;
        RECT 72.450 3311.390 82.110 3311.400 ;
        RECT 84.040 3311.390 85.880 3311.400 ;
        RECT 69.980 3310.940 85.880 3311.390 ;
        RECT 87.830 3311.290 88.180 3323.990 ;
        RECT 89.630 3317.270 90.030 3325.870 ;
        RECT 92.580 3323.170 94.580 3326.070 ;
        RECT 88.830 3316.870 90.030 3317.270 ;
        RECT 98.185 3313.670 98.780 3331.120 ;
        RECT 109.180 3319.520 109.660 3321.330 ;
        RECT 110.380 3320.870 110.780 3332.070 ;
        RECT 111.880 3332.070 116.880 3332.470 ;
        RECT 111.880 3321.320 112.380 3332.070 ;
        RECT 115.780 3330.070 116.180 3330.570 ;
        RECT 119.530 3330.120 119.930 3330.620 ;
        RECT 120.230 3330.420 120.630 3330.570 ;
        RECT 122.030 3330.420 122.430 3330.570 ;
        RECT 120.230 3329.920 122.430 3330.420 ;
        RECT 125.030 3330.120 125.430 3330.620 ;
        RECT 125.730 3330.470 126.130 3330.570 ;
        RECT 127.530 3330.470 127.930 3330.570 ;
        RECT 120.230 3329.770 120.630 3329.920 ;
        RECT 122.030 3329.770 122.430 3329.920 ;
        RECT 125.730 3329.920 127.930 3330.470 ;
        RECT 125.730 3329.770 126.130 3329.920 ;
        RECT 127.530 3329.770 127.930 3329.920 ;
        RECT 117.380 3326.870 117.780 3329.770 ;
        RECT 121.130 3328.870 123.330 3329.370 ;
        RECT 121.130 3328.770 121.530 3328.870 ;
        RECT 122.930 3328.770 123.330 3328.870 ;
        RECT 126.630 3328.770 128.830 3329.370 ;
        RECT 130.530 3326.870 130.930 3330.570 ;
        RECT 137.830 3330.320 138.330 3333.220 ;
        RECT 139.980 3331.470 144.430 3331.970 ;
        RECT 137.830 3329.820 138.830 3330.320 ;
        RECT 131.230 3326.870 131.630 3329.720 ;
        RECT 117.380 3326.470 131.630 3326.870 ;
        RECT 137.830 3325.920 138.330 3329.820 ;
        RECT 139.980 3327.720 140.480 3331.470 ;
        RECT 145.030 3330.970 145.530 3334.420 ;
        RECT 145.970 3332.040 157.930 3332.520 ;
        RECT 148.230 3332.020 150.680 3332.040 ;
        RECT 151.140 3331.500 151.430 3331.545 ;
        RECT 153.240 3331.500 153.530 3331.545 ;
        RECT 154.810 3331.500 155.100 3331.545 ;
        RECT 151.140 3331.360 155.100 3331.500 ;
        RECT 151.140 3331.315 151.430 3331.360 ;
        RECT 153.240 3331.315 153.530 3331.360 ;
        RECT 154.810 3331.315 155.100 3331.360 ;
        RECT 151.535 3331.160 151.825 3331.205 ;
        RECT 152.725 3331.160 153.015 3331.205 ;
        RECT 155.245 3331.160 155.535 3331.205 ;
        RECT 151.535 3331.020 155.535 3331.160 ;
        RECT 151.535 3330.975 151.825 3331.020 ;
        RECT 152.725 3330.975 153.015 3331.020 ;
        RECT 155.245 3330.975 155.535 3331.020 ;
        RECT 143.280 3330.670 146.480 3330.970 ;
        RECT 143.280 3328.970 143.580 3330.670 ;
        RECT 146.080 3330.570 146.480 3330.670 ;
        RECT 151.830 3330.420 152.330 3330.770 ;
        RECT 144.030 3329.820 144.430 3330.320 ;
        RECT 149.180 3330.070 152.330 3330.420 ;
        RECT 149.180 3329.870 149.730 3330.070 ;
        RECT 157.480 3329.970 165.680 3330.470 ;
        RECT 145.970 3329.670 148.270 3329.800 ;
        RECT 150.570 3329.720 157.930 3329.800 ;
        RECT 150.570 3329.670 162.680 3329.720 ;
        RECT 145.970 3329.320 162.680 3329.670 ;
        RECT 143.280 3328.670 147.230 3328.970 ;
        RECT 143.030 3327.870 146.530 3328.320 ;
        RECT 143.030 3327.720 143.430 3327.870 ;
        RECT 143.770 3327.840 146.530 3327.870 ;
        RECT 139.980 3327.220 143.430 3327.720 ;
        RECT 146.930 3326.620 147.230 3328.670 ;
        RECT 158.830 3328.320 159.230 3328.820 ;
        RECT 147.680 3327.870 159.230 3328.320 ;
        RECT 149.170 3327.840 159.230 3327.870 ;
        RECT 158.830 3327.820 159.230 3327.840 ;
        RECT 159.580 3327.670 160.080 3328.820 ;
        RECT 156.030 3327.420 160.080 3327.670 ;
        RECT 149.740 3327.300 150.030 3327.345 ;
        RECT 151.840 3327.300 152.130 3327.345 ;
        RECT 153.410 3327.300 153.700 3327.345 ;
        RECT 149.740 3327.160 153.700 3327.300 ;
        RECT 149.740 3327.115 150.030 3327.160 ;
        RECT 151.840 3327.115 152.130 3327.160 ;
        RECT 153.410 3327.115 153.700 3327.160 ;
        RECT 149.230 3326.620 149.630 3326.970 ;
        RECT 150.135 3326.960 150.425 3327.005 ;
        RECT 151.325 3326.960 151.615 3327.005 ;
        RECT 153.845 3326.960 154.135 3327.005 ;
        RECT 150.135 3326.820 154.135 3326.960 ;
        RECT 150.135 3326.775 150.425 3326.820 ;
        RECT 151.325 3326.775 151.615 3326.820 ;
        RECT 153.845 3326.775 154.135 3326.820 ;
        RECT 146.930 3326.320 149.630 3326.620 ;
        RECT 150.530 3326.070 150.930 3326.670 ;
        RECT 137.830 3325.570 143.430 3325.920 ;
        RECT 148.180 3325.820 150.930 3326.070 ;
        RECT 156.030 3326.620 156.480 3327.420 ;
        RECT 159.180 3326.870 159.680 3327.270 ;
        RECT 156.030 3325.870 156.530 3326.620 ;
        RECT 143.770 3325.570 146.530 3325.600 ;
        RECT 137.830 3325.420 146.530 3325.570 ;
        RECT 119.630 3324.120 125.030 3324.620 ;
        RECT 116.130 3323.070 116.530 3323.570 ;
        RECT 116.830 3323.370 117.230 3323.520 ;
        RECT 118.630 3323.370 119.030 3323.520 ;
        RECT 116.830 3322.870 119.030 3323.370 ;
        RECT 116.830 3322.720 117.230 3322.870 ;
        RECT 118.630 3322.720 119.030 3322.870 ;
        RECT 111.900 3319.520 112.380 3321.320 ;
        RECT 116.830 3320.170 117.230 3320.320 ;
        RECT 118.630 3320.170 119.030 3320.320 ;
        RECT 116.830 3319.670 119.030 3320.170 ;
        RECT 116.830 3319.520 117.230 3319.670 ;
        RECT 118.630 3319.520 119.030 3319.670 ;
        RECT 109.180 3319.170 109.680 3319.520 ;
        RECT 111.880 3319.270 112.380 3319.520 ;
        RECT 109.180 3318.770 110.180 3319.170 ;
        RECT 111.080 3318.870 112.380 3319.270 ;
        RECT 119.630 3319.120 120.130 3324.120 ;
        RECT 109.180 3318.020 109.680 3318.770 ;
        RECT 111.880 3318.020 112.380 3318.870 ;
        RECT 117.230 3318.620 120.130 3319.120 ;
        RECT 120.930 3319.420 121.330 3323.420 ;
        RECT 121.630 3323.170 122.030 3323.370 ;
        RECT 123.430 3323.170 123.830 3323.370 ;
        RECT 121.630 3322.670 123.830 3323.170 ;
        RECT 121.630 3322.520 122.030 3322.670 ;
        RECT 123.430 3322.520 123.830 3322.670 ;
        RECT 124.530 3320.970 125.030 3324.120 ;
        RECT 125.480 3322.870 125.880 3323.370 ;
        RECT 127.280 3322.870 127.680 3323.370 ;
        RECT 129.980 3322.920 130.380 3323.420 ;
        RECT 130.680 3323.320 131.080 3323.470 ;
        RECT 132.480 3323.320 132.880 3323.470 ;
        RECT 125.480 3322.370 127.680 3322.870 ;
        RECT 130.680 3322.820 132.880 3323.320 ;
        RECT 130.680 3322.670 131.080 3322.820 ;
        RECT 132.480 3322.670 132.880 3322.820 ;
        RECT 125.480 3322.220 125.880 3322.370 ;
        RECT 127.280 3322.220 127.680 3322.370 ;
        RECT 122.030 3320.470 123.430 3320.970 ;
        RECT 124.530 3320.470 127.280 3320.970 ;
        RECT 127.980 3319.420 128.380 3321.820 ;
        RECT 130.680 3320.120 131.080 3320.270 ;
        RECT 132.480 3320.120 132.880 3320.270 ;
        RECT 130.680 3319.620 132.880 3320.120 ;
        RECT 130.680 3319.470 131.080 3319.620 ;
        RECT 132.480 3319.470 132.880 3319.620 ;
        RECT 120.930 3319.020 128.380 3319.420 ;
        RECT 109.180 3316.650 109.660 3318.020 ;
        RECT 110.780 3317.170 111.630 3317.520 ;
        RECT 98.180 3313.070 98.780 3313.670 ;
        RECT 109.230 3313.470 109.630 3316.650 ;
        RECT 110.780 3315.520 111.280 3317.170 ;
        RECT 111.900 3316.650 112.380 3318.020 ;
        RECT 117.530 3317.370 118.330 3318.070 ;
        RECT 116.480 3313.470 116.880 3315.870 ;
        RECT 117.730 3314.170 118.130 3317.370 ;
        RECT 120.930 3315.470 121.330 3319.020 ;
        RECT 131.080 3318.570 132.880 3319.070 ;
        RECT 132.480 3316.620 132.880 3318.570 ;
        RECT 137.830 3314.220 138.330 3325.420 ;
        RECT 143.030 3325.120 146.530 3325.420 ;
        RECT 139.980 3319.770 144.430 3320.270 ;
        RECT 139.980 3316.020 140.480 3319.770 ;
        RECT 144.930 3319.270 145.430 3323.570 ;
        RECT 148.180 3322.570 148.680 3325.820 ;
        RECT 159.080 3325.720 159.580 3326.120 ;
        RECT 149.170 3325.570 158.830 3325.600 ;
        RECT 162.230 3325.570 162.680 3329.320 ;
        RECT 149.170 3325.120 162.680 3325.570 ;
        RECT 165.180 3322.570 165.680 3329.970 ;
        RECT 148.180 3322.070 165.680 3322.570 ;
        RECT 145.970 3320.340 157.930 3320.820 ;
        RECT 148.230 3320.320 150.680 3320.340 ;
        RECT 151.140 3319.800 151.430 3319.845 ;
        RECT 153.240 3319.800 153.530 3319.845 ;
        RECT 154.810 3319.800 155.100 3319.845 ;
        RECT 151.140 3319.660 155.100 3319.800 ;
        RECT 151.140 3319.615 151.430 3319.660 ;
        RECT 153.240 3319.615 153.530 3319.660 ;
        RECT 154.810 3319.615 155.100 3319.660 ;
        RECT 151.535 3319.460 151.825 3319.505 ;
        RECT 152.725 3319.460 153.015 3319.505 ;
        RECT 155.245 3319.460 155.535 3319.505 ;
        RECT 151.535 3319.320 155.535 3319.460 ;
        RECT 151.535 3319.275 151.825 3319.320 ;
        RECT 152.725 3319.275 153.015 3319.320 ;
        RECT 155.245 3319.275 155.535 3319.320 ;
        RECT 143.280 3318.970 146.480 3319.270 ;
        RECT 143.280 3317.270 143.580 3318.970 ;
        RECT 146.080 3318.870 146.480 3318.970 ;
        RECT 151.830 3318.720 152.330 3319.070 ;
        RECT 144.030 3318.120 144.430 3318.620 ;
        RECT 149.180 3318.370 152.330 3318.720 ;
        RECT 149.180 3318.170 149.730 3318.370 ;
        RECT 157.480 3318.270 165.680 3318.770 ;
        RECT 145.970 3317.970 148.270 3318.100 ;
        RECT 150.570 3318.020 157.930 3318.100 ;
        RECT 150.570 3317.970 162.680 3318.020 ;
        RECT 145.970 3317.620 162.680 3317.970 ;
        RECT 143.280 3316.970 147.230 3317.270 ;
        RECT 143.030 3316.170 146.530 3316.620 ;
        RECT 143.030 3316.020 143.430 3316.170 ;
        RECT 143.770 3316.140 146.530 3316.170 ;
        RECT 139.980 3315.520 143.430 3316.020 ;
        RECT 146.930 3314.920 147.230 3316.970 ;
        RECT 158.830 3316.620 159.230 3317.120 ;
        RECT 147.680 3316.170 159.230 3316.620 ;
        RECT 149.170 3316.140 159.230 3316.170 ;
        RECT 158.830 3316.120 159.230 3316.140 ;
        RECT 159.580 3316.770 160.630 3317.270 ;
        RECT 159.580 3315.970 160.080 3316.770 ;
        RECT 156.030 3315.720 160.080 3315.970 ;
        RECT 149.740 3315.600 150.030 3315.645 ;
        RECT 151.840 3315.600 152.130 3315.645 ;
        RECT 153.410 3315.600 153.700 3315.645 ;
        RECT 149.740 3315.460 153.700 3315.600 ;
        RECT 149.740 3315.415 150.030 3315.460 ;
        RECT 151.840 3315.415 152.130 3315.460 ;
        RECT 153.410 3315.415 153.700 3315.460 ;
        RECT 149.230 3314.920 149.630 3315.270 ;
        RECT 150.135 3315.260 150.425 3315.305 ;
        RECT 151.325 3315.260 151.615 3315.305 ;
        RECT 153.845 3315.260 154.135 3315.305 ;
        RECT 150.135 3315.120 154.135 3315.260 ;
        RECT 150.135 3315.075 150.425 3315.120 ;
        RECT 151.325 3315.075 151.615 3315.120 ;
        RECT 153.845 3315.075 154.135 3315.120 ;
        RECT 146.930 3314.620 149.630 3314.920 ;
        RECT 150.530 3314.370 150.930 3314.970 ;
        RECT 117.730 3314.100 119.180 3314.170 ;
        RECT 117.730 3313.850 121.145 3314.100 ;
        RECT 129.595 3313.850 131.700 3314.100 ;
        RECT 137.830 3313.870 143.430 3314.220 ;
        RECT 148.180 3314.120 150.930 3314.370 ;
        RECT 156.030 3314.920 156.480 3315.720 ;
        RECT 159.180 3315.170 159.680 3315.570 ;
        RECT 156.030 3314.170 156.530 3314.920 ;
        RECT 143.770 3313.870 146.530 3313.900 ;
        RECT 117.730 3313.770 119.180 3313.850 ;
        RECT 137.830 3313.720 146.530 3313.870 ;
        RECT 109.230 3313.070 118.680 3313.470 ;
        RECT 97.580 3312.470 98.780 3313.070 ;
        RECT 87.430 3310.940 88.180 3311.290 ;
        RECT 69.980 3310.920 71.980 3310.940 ;
        RECT 72.450 3310.920 83.080 3310.940 ;
        RECT 84.040 3310.920 85.880 3310.940 ;
        RECT 77.430 3310.370 79.430 3310.920 ;
        RECT 68.980 3308.920 70.180 3310.020 ;
        RECT 68.980 3307.770 70.980 3308.920 ;
        RECT 118.180 3308.820 118.680 3313.070 ;
        RECT 137.830 3308.820 138.330 3313.720 ;
        RECT 143.030 3313.420 146.530 3313.720 ;
        RECT 148.180 3310.870 148.680 3314.120 ;
        RECT 159.080 3314.020 159.580 3314.420 ;
        RECT 149.170 3313.870 158.830 3313.900 ;
        RECT 162.230 3313.870 162.680 3317.620 ;
        RECT 149.170 3313.420 162.680 3313.870 ;
        RECT 165.180 3310.870 165.680 3318.270 ;
        RECT 148.180 3310.370 165.680 3310.870 ;
        RECT 170.730 3308.820 171.230 3347.870 ;
        RECT 118.180 3308.320 171.230 3308.820 ;
        RECT 163.530 3306.520 164.030 3306.920 ;
        RECT 66.980 3306.120 164.030 3306.520 ;
      LAYER met2 ;
        RECT 74.630 3396.570 76.630 3397.670 ;
        RECT 94.280 3396.570 96.280 3397.670 ;
        RECT 133.380 3396.570 135.380 3397.720 ;
        RECT 157.530 3396.570 159.530 3397.670 ;
        RECT 151.580 3378.120 153.130 3380.120 ;
        RECT 70.780 3360.170 72.780 3362.170 ;
        RECT 76.580 3360.170 78.580 3362.170 ;
        RECT 82.630 3360.170 84.630 3362.170 ;
        RECT 76.130 3353.590 76.630 3354.140 ;
        RECT 76.130 3352.440 76.480 3353.590 ;
        RECT 72.980 3352.090 76.480 3352.440 ;
        RECT 70.130 3349.340 70.580 3349.390 ;
        RECT 72.980 3349.340 73.330 3352.090 ;
        RECT 70.130 3348.990 73.330 3349.340 ;
        RECT 70.130 3348.940 70.580 3348.990 ;
        RECT 72.980 3347.040 73.330 3348.990 ;
        RECT 72.980 3346.690 78.380 3347.040 ;
        RECT 78.030 3345.090 78.380 3346.690 ;
        RECT 78.030 3344.590 78.530 3345.090 ;
        RECT 89.980 3339.470 91.980 3341.220 ;
        RECT 115.280 3337.620 115.780 3349.820 ;
        RECT 170.730 3342.920 172.130 3344.920 ;
        RECT 143.980 3337.620 145.280 3338.920 ;
        RECT 115.280 3337.170 145.280 3337.620 ;
        RECT 66.580 3333.670 68.580 3335.670 ;
        RECT 69.330 3332.620 70.330 3335.670 ;
        RECT 41.280 3331.620 70.330 3332.620 ;
        RECT 115.280 3332.070 115.780 3337.170 ;
        RECT 143.980 3336.920 145.280 3337.170 ;
        RECT 41.280 3230.350 43.280 3331.620 ;
        RECT 70.780 3327.270 72.780 3329.270 ;
        RECT 79.430 3327.270 81.430 3329.270 ;
        RECT 88.630 3327.270 90.630 3329.270 ;
        RECT 159.580 3328.320 164.230 3328.820 ;
        RECT 92.180 3326.070 94.180 3326.120 ;
        RECT 76.130 3321.940 76.630 3322.490 ;
        RECT 68.380 3320.020 70.780 3321.320 ;
        RECT 76.130 3320.790 76.480 3321.940 ;
        RECT 72.980 3320.440 76.480 3320.790 ;
        RECT 70.130 3317.690 70.580 3317.740 ;
        RECT 72.980 3317.690 73.330 3320.440 ;
        RECT 70.130 3317.340 73.330 3317.690 ;
        RECT 64.180 3313.420 65.180 3317.320 ;
        RECT 70.130 3317.290 70.580 3317.340 ;
        RECT 72.980 3315.390 73.330 3317.340 ;
        RECT 72.980 3315.040 78.380 3315.390 ;
        RECT 78.030 3313.440 78.380 3315.040 ;
        RECT 64.180 3312.420 68.280 3313.420 ;
        RECT 78.030 3312.940 78.530 3313.440 ;
        RECT 66.280 3236.120 68.280 3312.420 ;
        RECT 77.430 3309.820 79.430 3310.920 ;
        RECT 68.980 3307.770 70.980 3308.870 ;
        RECT 66.280 3234.120 74.230 3236.120 ;
        RECT 72.230 3230.350 74.230 3234.120 ;
        RECT 92.180 3230.830 94.580 3326.070 ;
        RECT 163.730 3323.570 164.230 3328.320 ;
        RECT 144.930 3323.070 164.230 3323.570 ;
        RECT 170.730 3319.920 171.980 3321.920 ;
        RECT 128.180 3307.620 130.130 3308.820 ;
        RECT 158.530 3307.620 160.480 3308.820 ;
        RECT 41.150 3223.450 43.450 3230.350 ;
        RECT 71.940 3223.450 74.700 3230.350 ;
        RECT 92.180 3223.470 94.940 3230.830 ;
      LAYER met3 ;
        RECT 33.530 3413.320 202.980 3416.420 ;
        RECT 57.380 3403.120 178.930 3406.120 ;
        RECT 74.630 3396.970 76.630 3398.470 ;
        RECT 94.280 3396.970 96.280 3398.470 ;
        RECT 133.380 3396.970 135.380 3398.470 ;
        RECT 157.530 3396.970 159.530 3398.370 ;
        RECT 151.580 3378.120 178.930 3380.120 ;
        RECT 33.530 3360.170 84.630 3362.170 ;
        RECT 170.730 3342.920 178.930 3344.920 ;
        RECT 57.530 3339.220 91.980 3341.220 ;
        RECT 143.980 3336.970 202.980 3338.920 ;
        RECT 143.980 3336.920 197.930 3336.970 ;
        RECT 33.530 3333.670 68.580 3335.670 ;
        RECT 61.730 3327.270 90.630 3329.270 ;
        RECT 61.730 3325.320 63.830 3327.270 ;
        RECT 60.930 3325.270 63.830 3325.320 ;
        RECT 57.530 3323.270 63.830 3325.270 ;
        RECT 57.530 3320.020 70.780 3321.470 ;
        RECT 57.530 3319.470 60.180 3320.020 ;
        RECT 170.730 3319.920 178.930 3321.920 ;
        RECT 77.430 3309.220 79.430 3310.420 ;
        RECT 68.980 3307.120 70.980 3308.420 ;
        RECT 128.180 3307.070 130.130 3308.320 ;
        RECT 158.530 3306.920 160.480 3308.320 ;
        RECT 57.380 3261.020 178.930 3264.120 ;
        RECT 33.530 3239.220 202.980 3242.220 ;
      LAYER met4 ;
        RECT 33.530 3239.220 36.630 3416.420 ;
        RECT 57.380 3261.020 60.380 3406.120 ;
        RECT 74.630 3396.570 76.630 3416.420 ;
        RECT 94.280 3396.570 96.280 3416.420 ;
        RECT 133.380 3396.570 135.380 3416.420 ;
        RECT 157.530 3396.570 159.530 3416.420 ;
        RECT 199.980 3416.120 202.980 3416.420 ;
        RECT 175.780 3405.920 178.930 3406.120 ;
        RECT 68.980 3239.220 70.980 3308.870 ;
        RECT 77.430 3239.270 79.430 3310.920 ;
        RECT 128.180 3261.045 130.130 3308.870 ;
        RECT 158.530 3261.045 160.480 3308.820 ;
        RECT 175.760 3261.120 178.930 3405.920 ;
        RECT 175.780 3261.020 178.930 3261.120 ;
        RECT 199.960 3239.240 202.980 3416.120 ;
        RECT 199.980 3239.220 202.980 3239.240 ;
  END
END user_project_wrapper
END LIBRARY

