magic
tech sky130A
timestamp 1724038531
<< nwell >>
rect -30 1015 -10 1035
rect -30 975 -10 995
rect 780 815 800 835
rect 810 795 825 815
rect 830 525 890 1105
rect 920 1015 940 1035
rect 1400 1015 1420 1035
rect 1840 995 1940 1105
rect 1945 1015 1965 1035
rect 920 975 940 995
rect 1400 975 1420 995
rect 1840 975 1935 995
rect 1945 975 1965 995
rect 1335 955 1355 965
rect 1325 935 1355 955
rect 1335 920 1355 935
rect 1840 940 1940 975
rect 1840 915 1935 940
rect 1850 865 1925 915
rect 1805 655 1825 675
rect 1840 525 1940 865
rect 2730 855 2745 865
rect 2755 855 2775 875
rect 2730 845 2755 855
<< pwell >>
rect -60 -20 2805 460
rect -40 -40 0 -20
<< pmos >>
rect 2730 845 2745 865
<< ndiff >>
rect 2745 430 2785 440
<< pdiff >>
rect 1335 955 1355 965
rect 1345 935 1355 955
rect 1335 920 1355 935
rect 2745 845 2755 855
<< ndiffc >>
rect 1805 330 1825 350
rect 2755 330 2775 350
rect -30 90 -10 110
rect 920 90 940 110
rect 1400 90 1420 110
rect 1945 90 1965 110
rect -30 50 -10 70
rect 920 50 940 70
rect 1400 50 1420 70
rect 1945 50 1965 70
<< pdiffc >>
rect -30 1015 -10 1035
rect 920 1015 940 1035
rect 1400 1015 1420 1035
rect 1945 1015 1965 1035
rect -30 975 -10 995
rect 920 975 940 995
rect 1400 975 1420 995
rect 1945 975 1965 995
rect 1325 935 1345 955
rect 2755 855 2775 875
rect 780 815 800 835
rect 1805 655 1825 675
<< psubdiff >>
rect 840 150 880 165
rect 840 130 850 150
rect 870 130 880 150
rect 840 110 880 130
rect 1865 150 1905 165
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 1865 110 1905 130
rect 840 90 850 110
rect 870 90 880 110
rect 1865 90 1875 110
rect 1895 90 1905 110
rect 840 70 880 90
rect 1865 70 1905 90
rect 840 50 850 70
rect 870 50 880 70
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 840 35 880 50
rect 1865 35 1905 50
<< nsubdiff >>
rect 840 1035 880 1050
rect 1865 1045 1905 1060
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 840 995 880 1015
rect 1865 1005 1905 1025
rect 840 975 850 995
rect 870 975 880 995
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 840 955 880 975
rect 1865 965 1905 985
rect 840 935 850 955
rect 870 935 880 955
rect 840 920 880 935
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 1865 930 1905 945
<< psubdiffcont >>
rect 850 130 870 150
rect 1875 130 1895 150
rect 850 90 870 110
rect 1875 90 1895 110
rect 850 50 870 70
rect 1875 50 1895 70
<< nsubdiffcont >>
rect 850 1015 870 1035
rect 1875 1025 1895 1045
rect 850 975 870 995
rect 1875 985 1895 1005
rect 850 935 870 955
rect 1875 945 1895 965
<< poly >>
rect 170 505 190 515
rect 365 470 405 515
rect 2340 470 2380 515
rect 2735 470 2745 515
<< polycont >>
rect 10 480 30 500
rect 50 480 70 500
rect 90 480 110 500
rect 130 480 150 500
rect 170 480 190 500
rect 210 480 230 500
rect 250 480 270 500
rect 290 480 310 500
rect 330 480 350 500
rect 420 480 440 500
rect 460 480 480 500
rect 500 480 520 500
rect 540 480 560 500
rect 580 480 600 500
rect 620 480 640 500
rect 660 480 680 500
rect 700 480 720 500
rect 740 480 760 500
rect 960 480 980 500
rect 1000 480 1020 500
rect 1040 480 1060 500
rect 1080 480 1100 500
rect 1120 480 1140 500
rect 1160 480 1180 500
rect 1200 480 1220 500
rect 1240 480 1260 500
rect 1280 480 1300 500
rect 1440 480 1460 500
rect 1480 480 1500 500
rect 1520 480 1540 500
rect 1560 480 1580 500
rect 1600 480 1620 500
rect 1640 480 1660 500
rect 1680 480 1700 500
rect 1720 480 1740 500
rect 1760 480 1780 500
rect 1985 480 2005 500
rect 2025 480 2045 500
rect 2065 480 2085 500
rect 2105 480 2125 500
rect 2145 480 2165 500
rect 2185 480 2205 500
rect 2225 480 2245 500
rect 2265 480 2285 500
rect 2305 480 2325 500
rect 2390 480 2410 500
rect 2430 480 2450 500
rect 2470 480 2490 500
rect 2510 480 2530 500
rect 2550 480 2570 500
rect 2590 480 2610 500
rect 2630 480 2650 500
rect 2670 480 2690 500
rect 2710 480 2730 500
<< locali >>
rect 840 1035 880 1050
rect 1865 1045 1905 1060
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 840 995 880 1015
rect 1865 1005 1905 1025
rect 840 975 850 995
rect 870 975 880 995
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 2340 995 2380 1045
rect 840 955 880 975
rect 1865 965 1905 985
rect 1335 955 1355 965
rect 840 935 850 955
rect 870 935 880 955
rect 1345 935 1355 955
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 2340 960 2380 975
rect 840 920 880 935
rect 1335 920 1355 935
rect 1865 930 1905 945
rect 2375 940 2380 960
rect 2340 545 2380 865
rect 2745 845 2755 855
rect 2755 575 2775 595
rect 0 500 770 515
rect 0 480 10 500
rect 30 480 50 500
rect 70 480 90 500
rect 110 480 130 500
rect 150 480 170 500
rect 190 480 210 500
rect 230 480 250 500
rect 270 480 290 500
rect 310 480 330 500
rect 350 480 420 500
rect 440 480 460 500
rect 480 480 500 500
rect 520 480 540 500
rect 560 480 580 500
rect 600 480 620 500
rect 640 480 660 500
rect 680 480 700 500
rect 720 480 740 500
rect 760 480 770 500
rect 0 470 770 480
rect 790 440 810 545
rect 950 500 1315 515
rect 950 480 960 500
rect 980 480 1000 500
rect 1020 480 1040 500
rect 1060 480 1080 500
rect 1100 480 1120 500
rect 1140 480 1160 500
rect 1180 480 1200 500
rect 1220 480 1240 500
rect 1260 480 1280 500
rect 1300 480 1315 500
rect 950 470 1315 480
rect 1335 440 1355 545
rect 1430 500 1795 515
rect 1430 480 1440 500
rect 1460 480 1480 500
rect 1500 480 1520 500
rect 1540 480 1560 500
rect 1580 480 1600 500
rect 1620 480 1640 500
rect 1660 480 1680 500
rect 1700 480 1720 500
rect 1740 480 1760 500
rect 1780 480 1795 500
rect 1430 470 1795 480
rect 1815 440 1835 545
rect 1975 500 2745 515
rect 1975 480 1985 500
rect 2005 480 2025 500
rect 2045 480 2065 500
rect 2085 480 2105 500
rect 2125 480 2145 500
rect 2165 480 2185 500
rect 2205 480 2225 500
rect 2245 480 2265 500
rect 2285 480 2305 500
rect 2325 480 2390 500
rect 2410 480 2430 500
rect 2450 480 2470 500
rect 2490 480 2510 500
rect 2530 480 2550 500
rect 2570 480 2590 500
rect 2610 480 2630 500
rect 2650 480 2670 500
rect 2690 480 2710 500
rect 2730 480 2745 500
rect 1975 470 2745 480
rect 2765 440 2785 545
rect 2745 430 2785 440
rect 840 150 880 165
rect 1865 150 1905 165
rect 840 130 850 150
rect 870 130 880 150
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 840 110 880 130
rect 1865 110 1905 130
rect 840 90 850 110
rect 870 90 880 110
rect 1865 90 1875 110
rect 1895 90 1905 110
rect 840 70 880 90
rect 1865 70 1905 90
rect 840 50 850 70
rect 870 50 880 70
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 840 35 880 50
rect 1865 35 1905 50
<< viali >>
rect -30 1015 -10 1035
rect 850 1015 870 1035
rect 920 1015 940 1035
rect 1400 1015 1420 1035
rect 1875 1025 1895 1045
rect 1945 1015 1965 1035
rect -30 975 -10 995
rect 850 975 870 995
rect 920 975 940 995
rect 1400 975 1420 995
rect 1875 985 1895 1005
rect 1945 975 1965 995
rect -30 935 -10 955
rect 850 935 870 955
rect 920 935 940 955
rect 1325 935 1345 955
rect 1400 935 1420 955
rect 1875 945 1895 965
rect 1945 935 1965 955
rect 2755 935 2775 955
rect 1325 855 1345 875
rect 780 815 800 835
rect 1805 815 1825 835
rect 780 775 800 795
rect 1805 775 1825 795
rect 780 655 800 675
rect 1325 655 1345 675
rect 1805 655 1825 675
rect 780 575 800 595
rect 1325 575 1345 595
rect 1805 575 1825 595
rect 2755 855 2775 875
rect 10 480 30 500
rect 90 480 110 500
rect 170 480 190 500
rect 250 480 270 500
rect 330 480 350 500
rect 420 480 440 500
rect 500 480 520 500
rect 580 480 600 500
rect 660 480 680 500
rect 740 480 760 500
rect 960 480 980 500
rect 1040 480 1060 500
rect 1120 480 1140 500
rect 1200 480 1220 500
rect 1280 480 1300 500
rect 1440 480 1460 500
rect 1520 480 1540 500
rect 1600 480 1620 500
rect 1680 480 1700 500
rect 1760 480 1780 500
rect 1985 480 2005 500
rect 2065 480 2085 500
rect 2145 480 2165 500
rect 2225 480 2245 500
rect 2305 480 2325 500
rect 2390 480 2410 500
rect 2470 480 2490 500
rect 2550 480 2570 500
rect 2630 480 2650 500
rect 2710 480 2730 500
rect 780 410 800 430
rect 1325 410 1345 430
rect 1805 410 1825 430
rect 2755 410 2775 430
rect 780 330 800 350
rect 1325 330 1345 350
rect 1805 330 1825 350
rect 2755 330 2775 350
rect 2755 250 2775 270
rect -30 130 -10 150
rect 850 130 870 150
rect 920 130 940 150
rect 1400 130 1420 150
rect 1875 130 1895 150
rect 1945 130 1965 150
rect -30 90 -10 110
rect 850 90 870 110
rect 920 90 940 110
rect 1400 90 1420 110
rect 1875 90 1895 110
rect 1945 90 1965 110
rect -30 50 -10 70
rect 850 50 870 70
rect 920 50 940 70
rect 1400 50 1420 70
rect 1875 50 1895 70
rect 1945 50 1965 70
<< metal1 >>
rect -40 1035 0 1125
rect -40 1015 -30 1035
rect -10 1015 0 1035
rect -40 995 0 1015
rect -40 975 -30 995
rect -10 975 0 995
rect -40 955 0 975
rect -40 935 -30 955
rect -10 935 0 955
rect -40 925 0 935
rect 840 1035 880 1125
rect 840 1015 850 1035
rect 870 1015 880 1035
rect 840 995 880 1015
rect 840 975 850 995
rect 870 975 880 995
rect 840 955 880 975
rect 840 935 850 955
rect 870 935 880 955
rect 840 920 880 935
rect 910 1035 950 1125
rect 910 1015 920 1035
rect 940 1015 950 1035
rect 910 995 950 1015
rect 910 975 920 995
rect 940 975 950 995
rect 910 955 950 975
rect 1390 1035 1430 1125
rect 1390 1015 1400 1035
rect 1420 1015 1430 1035
rect 1390 995 1430 1015
rect 1390 975 1400 995
rect 1420 975 1430 995
rect 910 935 920 955
rect 940 935 950 955
rect 910 925 950 935
rect 1315 955 1355 965
rect 1315 935 1325 955
rect 1345 935 1355 955
rect 1315 895 1355 935
rect 1390 955 1430 975
rect 1390 935 1400 955
rect 1420 935 1430 955
rect 1390 925 1430 935
rect 1865 1045 1905 1125
rect 1865 1025 1875 1045
rect 1895 1025 1905 1045
rect 1865 1005 1905 1025
rect 1865 985 1875 1005
rect 1895 985 1905 1005
rect 1865 965 1905 985
rect 1865 945 1875 965
rect 1895 945 1905 965
rect 1865 930 1905 945
rect 1935 1035 1975 1125
rect 1935 1015 1945 1035
rect 1965 1015 1975 1035
rect 1935 995 1975 1015
rect 1935 975 1945 995
rect 1965 975 1975 995
rect 1935 955 1975 975
rect 1935 935 1945 955
rect 1965 935 1975 955
rect 1935 925 1975 935
rect 2745 955 2785 965
rect 2745 935 2755 955
rect 2775 935 2785 955
rect 2745 895 2785 935
rect 1315 875 2785 895
rect 1315 855 1325 875
rect 1345 855 2755 875
rect 2775 855 2785 875
rect 1315 845 2785 855
rect 770 835 810 845
rect 770 815 780 835
rect 800 815 810 835
rect 1795 835 1835 845
rect 1795 815 1805 835
rect 1825 815 1835 835
rect -60 765 190 815
rect 770 795 2805 815
rect 770 775 780 795
rect 800 775 1805 795
rect 1825 775 2805 795
rect 770 765 2805 775
rect 140 515 190 765
rect 770 675 810 685
rect 770 655 780 675
rect 800 655 810 675
rect 770 595 810 655
rect 770 575 780 595
rect 800 575 810 595
rect 770 545 810 575
rect 1315 675 1355 685
rect 1315 655 1325 675
rect 1345 655 1355 675
rect 1315 595 1355 655
rect 1315 575 1325 595
rect 1345 575 1355 595
rect 1315 545 1355 575
rect 1795 675 1835 685
rect 1795 655 1805 675
rect 1825 655 1835 675
rect 1795 595 1835 655
rect 1795 575 1805 595
rect 1825 575 1835 595
rect 1795 545 1835 575
rect 2745 545 2785 605
rect 790 515 810 545
rect 1335 515 1355 545
rect 0 500 770 515
rect 0 480 10 500
rect 30 480 90 500
rect 110 480 170 500
rect 190 480 250 500
rect 270 480 330 500
rect 350 480 420 500
rect 440 480 500 500
rect 520 480 580 500
rect 600 480 660 500
rect 680 480 740 500
rect 760 480 770 500
rect 0 470 770 480
rect 790 500 1315 515
rect 790 480 960 500
rect 980 480 1040 500
rect 1060 480 1120 500
rect 1140 480 1200 500
rect 1220 480 1280 500
rect 1300 480 1315 500
rect 790 470 1315 480
rect 1335 500 1795 515
rect 1335 480 1440 500
rect 1460 480 1520 500
rect 1540 480 1600 500
rect 1620 480 1680 500
rect 1700 480 1760 500
rect 1780 480 1795 500
rect 1335 470 1795 480
rect 790 440 810 470
rect 1335 440 1355 470
rect 1815 440 1835 545
rect 1975 500 2745 515
rect 1975 480 1985 500
rect 2005 480 2065 500
rect 2085 480 2145 500
rect 2165 480 2225 500
rect 2245 480 2305 500
rect 2325 480 2390 500
rect 2410 480 2470 500
rect 2490 480 2550 500
rect 2570 480 2630 500
rect 2650 480 2710 500
rect 2730 480 2745 500
rect 1975 470 2745 480
rect 770 430 810 440
rect 770 410 780 430
rect 800 410 810 430
rect 770 350 810 410
rect 770 330 780 350
rect 800 330 810 350
rect 770 320 810 330
rect 1315 430 1355 440
rect 1315 410 1325 430
rect 1345 410 1355 430
rect 1315 350 1355 410
rect 1315 330 1325 350
rect 1345 330 1355 350
rect 1315 320 1355 330
rect 1795 430 1835 440
rect 1795 410 1805 430
rect 1825 410 1835 430
rect 1795 350 1835 410
rect 1795 330 1805 350
rect 1825 330 1835 350
rect 1795 320 1835 330
rect 2105 290 2155 470
rect 2765 440 2785 545
rect -60 240 2155 290
rect 2745 430 2785 440
rect 2745 410 2755 430
rect 2775 410 2785 430
rect 2745 350 2785 410
rect 2745 330 2755 350
rect 2775 330 2785 350
rect 2745 290 2785 330
rect 2745 270 2805 290
rect 2745 250 2755 270
rect 2775 250 2805 270
rect 2745 240 2805 250
rect -40 150 0 160
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 -40 0 50
rect 840 150 880 165
rect 840 130 850 150
rect 870 130 880 150
rect 840 110 880 130
rect 840 90 850 110
rect 870 90 880 110
rect 840 70 880 90
rect 840 50 850 70
rect 870 50 880 70
rect 840 -40 880 50
rect 910 150 950 160
rect 910 130 920 150
rect 940 130 950 150
rect 910 110 950 130
rect 910 90 920 110
rect 940 90 950 110
rect 910 70 950 90
rect 910 50 920 70
rect 940 50 950 70
rect 910 -40 950 50
rect 1390 150 1430 160
rect 1390 130 1400 150
rect 1420 130 1430 150
rect 1390 110 1430 130
rect 1390 90 1400 110
rect 1420 90 1430 110
rect 1390 70 1430 90
rect 1390 50 1400 70
rect 1420 50 1430 70
rect 1390 -40 1430 50
rect 1865 150 1905 165
rect 1865 130 1875 150
rect 1895 130 1905 150
rect 1865 110 1905 130
rect 1865 90 1875 110
rect 1895 90 1905 110
rect 1865 70 1905 90
rect 1865 50 1875 70
rect 1895 50 1905 70
rect 1865 -40 1905 50
rect 1935 150 1975 160
rect 1935 130 1945 150
rect 1965 130 1975 150
rect 1935 110 1975 130
rect 1935 90 1945 110
rect 1965 90 1975 110
rect 1935 70 1975 90
rect 1935 50 1945 70
rect 1965 50 1975 70
rect 1935 -40 1975 50
use inv  inv_2
timestamp 1723457586
transform 1 0 950 0 1 545
box -60 -545 425 560
use inv  inv_3
timestamp 1723457586
transform 1 0 1430 0 1 545
box -60 -545 425 560
use main_inv_vco  main_inv_vco_0
timestamp 1724038090
transform 1 0 0 0 1 545
box -60 -545 830 560
use main_inv_vco  main_inv_vco_1
timestamp 1724038090
transform 1 0 1975 0 1 545
box -60 -545 830 560
<< labels >>
rlabel metal1 -60 805 -60 805 7 inp
port 1 w
rlabel metal1 -60 280 -60 280 7 inn
port 2 w
rlabel metal1 2805 805 2805 805 3 outp
port 3 e
rlabel metal1 2805 280 2805 280 3 outn
port 4 e
rlabel metal1 860 1125 860 1125 1 VCCA
port 5 n
rlabel metal1 1885 1125 1885 1125 1 VCCA
port 6 n
rlabel metal1 860 -40 860 -40 5 GND
port 7 s
rlabel metal1 1885 -40 1885 -40 5 GND
port 8 s
rlabel metal1 -20 1125 -20 1125 1 VPWR
port 9 n
rlabel metal1 930 1125 930 1125 1 VPWR
port 10 n
rlabel metal1 1410 1125 1410 1125 1 VPWR
port 11 n
rlabel metal1 1955 1125 1955 1125 1 VPWR
port 12 n
rlabel metal1 -20 -40 -20 -40 5 VGND
port 13 s
rlabel metal1 930 -40 930 -40 5 VGND
port 14 s
rlabel metal1 1410 -40 1410 -40 5 VGND
port 15 s
rlabel metal1 1955 -40 1955 -40 5 VGND
port 16 s
<< end >>
