* NGSPICE file created from dco.ext - technology: sky130A

.s

.subckt dco_freq clk clkDiv2 VNB VGND VPB VPWR
Xsky130_fd_sc_hd__buf_4_0 Q_N VGND VNB VPB VPWR Q_N_buf sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_4_0 clk VGND VNB VPB VPWR clkinv sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__dfxtp_1_0 clkinv Q_N_buf VGND VNB VPB VPWR D sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxbp_2_0 clk D VGND VNB VPB VPWR clkDiv2 Q_N sky130_fd_sc_hd__dfxbp_2
.ends


.subckt dco_aux_inv VPWR VCCA A Y GND VGND
X0 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1
X1 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=1
.ends

.subckt dco_main_inv VPWR VCCA Y GND VGND A
X0 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=1 M=2
X1 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=1 M=2
.ends

.subckt dco_cc_inv outp inp inn outn VCCA VGND VPWR GND
Xdco_aux_inv_0 VPWR VCCA outp outn GND VGND dco_aux_inv
Xdco_aux_inv_1 VPWR VCCA outn outp GND VGND dco_aux_inv
Xdco_main_inv_0 VPWR VCCA outp GND VGND inp dco_main_inv
Xdco_main_inv_1 VPWR VCCA outn GND VGND inn dco_main_inv
.ends

.subckt dco_ring_osc p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4] VGND p[0] VPWR
+ GND VCCA
Xdco_cc_inv_0 p[0] p[4] pn[4] pn[0] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_1 p[1] p[0] pn[0] pn[1] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_2 p[2] p[1] pn[1] pn[2] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_3 p[4] p[3] pn[3] pn[4] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_4 p[3] p[2] pn[2] pn[3] VCCA VGND VPWR GND dco_cc_inv
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_RSCMUS a_n35_n1272# a_n35_840# a_n165_n1402#
X0 a_n35_840# a_n35_n1272# a_n165_n1402# sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

.subckt dco_idac Dctrl Vbs1 Vbs2 Vbs3 Vbs4 Isup VCCD VCCA GND
Xsky130_fd_sc_hd__buf_2_0 Dctrl GND GND VCCD VCCD G_M7 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 G_M7 GND GND VCCD VCCD G_M5 sky130_fd_sc_hd__inv_2
Xsky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0 GND D_M7 GND sky130_fd_pr__res_xhigh_po_0p35_RSCMUS
X0 Isup G_M7 D1_M4 GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X1 B_M2 Vbs1 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X2 D1_M4 Vbs4 D1_M3 D1_M3 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X3 D_M7 G_M5 D1_M4 GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X4 Isup G_M5 D1_M4 D1_M4 sky130_fd_pr__pfet_01v8_hvt ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
X5 D1_M3 Vbs3 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X6 Isup Vbs2 B_M2 B_M2 sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X7 D1_M4 G_M7 D_M7 D1_M4 sky130_fd_pr__pfet_01v8_hvt ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.5 M=2
.ends


.subckt dco VCCD VCCA Dctrl ENB Vbs_12 Vbs_34 pha_DCO
Xdco_freq_0 pha_ro ro_div2 GND GND VCCD VCCD dco_freq
Xdco_freq_1 ro_div2 pha_DCO GND GND VCCD VCCD dco_freq
Xsky130_fd_sc_hd__buf_2_0 p_osc GND GND VCCD VCCD pha_ro sky130_fd_sc_hd__buf_2
Xdco_ring_osc_0 dco_ring_osc_0/p[1] dco_ring_osc_0/p[2] dco_ring_osc_0/p[3] p_osc
+ dco_ring_osc_0/pn[0] dco_ring_osc_0/pn[1] dco_ring_osc_0/pn[2] dco_ring_osc_0/pn[3]
+ dco_ring_osc_0/pn[4] GND dco_ring_osc_0/p[0] Isup GND Isup dco_ring_osc
Xdco_idac_0 Dctrl Vbs_12 Vbs_12 Vbs_34 Vbs_34 Isup VCCD VCCA GND dco_idac
Xsky130_fd_sc_hd__einvp_1_0 VCCD ENB GND GND VCCD VCCD dco_ring_osc_0/pn[4] sky130_fd_sc_hd__einvp_1
.ends

