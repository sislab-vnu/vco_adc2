* NGSPICE file created from count.ext - technology: sky130A


.subckt count UP SetB DOWN Dout_buf
Xsky130_fd_sc_hd__dfstp_1_0 UP_buf Q2N SetBi GND GND VCCD VCCD Q1 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfstp_1_1 sky130_fd_sc_hd__dfstp_1_1/CLK Q1_buf SetBi GND GND VCCD
+ VCCD Q2 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__buf_2_0 UP GND GND VCCD VCCD UP_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 SetB GND GND sky130_fd_sc_hd__inv_2_0/VPB VCCD SetBi sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_1 DOWN GND GND VCCD VCCD sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_1 Q2 GND GND VCCD VCCD Q2N sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_2 Dout GND GND VCCD VCCD Dout_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_3 Q1 GND GND VCCD VCCD Q1_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_1 Q1 Q2 GND GND VCCD VCCD Dout sky130_fd_sc_hd__xor2_1
.ends

