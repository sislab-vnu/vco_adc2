magic
tech sky130A
timestamp 1726545299
<< pwell >>
rect -130 -40 200 240
<< nmos >>
rect 0 0 50 200
rect 90 0 140 200
<< ndiff >>
rect -40 190 0 200
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 190 90 200
rect 50 170 60 190
rect 80 170 90 190
rect 50 150 90 170
rect 50 130 60 150
rect 80 130 90 150
rect 50 110 90 130
rect 50 90 60 110
rect 80 90 90 110
rect 50 70 90 90
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 190 180 200
rect 140 170 150 190
rect 170 170 180 190
rect 140 150 180 170
rect 140 130 150 150
rect 170 130 180 150
rect 140 110 180 130
rect 140 90 150 110
rect 170 90 180 110
rect 140 70 180 90
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
<< ndiffc >>
rect -30 170 -10 190
rect -30 130 -10 150
rect -30 90 -10 110
rect -30 50 -10 70
rect -30 10 -10 30
rect 60 170 80 190
rect 60 130 80 150
rect 60 90 80 110
rect 60 50 80 70
rect 60 10 80 30
rect 150 170 170 190
rect 150 130 170 150
rect 150 90 170 110
rect 150 50 170 70
rect 150 10 170 30
<< psubdiff >>
rect -110 190 -70 205
rect -110 170 -100 190
rect -80 170 -70 190
rect -110 155 -70 170
<< psubdiffcont >>
rect -100 170 -80 190
<< poly >>
rect 0 270 140 280
rect 0 250 40 270
rect 100 250 140 270
rect 0 240 140 250
rect 0 200 50 240
rect 90 200 140 240
rect 0 -40 50 0
rect 90 -40 140 0
<< polycont >>
rect 40 250 100 270
<< locali >>
rect 25 270 115 280
rect 25 250 40 270
rect 100 250 115 270
rect 25 240 115 250
rect -110 190 -70 205
rect -110 170 -100 190
rect -80 170 -70 190
rect -110 155 -70 170
rect -40 190 0 200
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 190 90 200
rect 50 170 60 190
rect 80 170 90 190
rect 50 150 90 170
rect 50 130 60 150
rect 80 130 90 150
rect 50 110 90 130
rect 50 90 60 110
rect 80 90 90 110
rect 50 70 90 90
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 190 180 200
rect 140 170 150 190
rect 170 170 180 190
rect 140 150 180 170
rect 140 130 150 150
rect 170 130 180 150
rect 140 110 180 130
rect 140 90 150 110
rect 170 90 180 110
rect 140 70 180 90
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
<< viali >>
rect 40 250 100 270
rect -100 170 -80 190
rect -30 170 -10 190
rect -30 130 -10 150
rect -30 50 -10 70
rect -30 10 -10 30
rect 150 170 170 190
rect 150 130 170 150
rect 150 50 170 70
rect 150 10 170 30
<< metal1 >>
rect 0 270 140 280
rect 0 250 40 270
rect 100 250 140 270
rect 0 240 140 250
rect -110 190 -70 205
rect -110 170 -100 190
rect -80 170 -70 190
rect -110 155 -70 170
rect -40 190 0 200
rect -40 170 -30 190
rect -10 185 0 190
rect 140 190 180 200
rect 140 185 150 190
rect -10 170 150 185
rect 170 170 180 190
rect -40 150 180 170
rect -40 130 -30 150
rect -10 135 150 150
rect -10 130 0 135
rect -40 120 0 130
rect 140 130 150 135
rect 170 130 180 150
rect 140 120 180 130
rect -40 70 0 80
rect -40 50 -30 70
rect -10 65 0 70
rect 140 70 180 80
rect 140 65 150 70
rect -10 50 150 65
rect 170 50 180 70
rect -40 30 180 50
rect -40 10 -30 30
rect -10 15 150 30
rect -10 10 0 15
rect -40 0 0 10
rect 140 10 150 15
rect 170 10 180 30
rect 140 0 180 10
<< labels >>
rlabel metal1 -90 205 -90 205 1 B
rlabel metal1 -20 200 -20 200 1 S
rlabel locali 70 0 70 0 5 D
rlabel metal1 70 280 70 280 1 G
<< end >>
