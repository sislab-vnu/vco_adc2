* Cell		: DCO design
* Written for	: NGSPICE
* Lib		:  Testbenchs
******************************************************

.lib /home/dkit/efabless/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc ../library/analog_lib_for_design.spice
.inc ../library/digital_lib.spice
*.option savecurrents
.global gnd vdd
.param mc_mm_switch=0
*---------- sub circuits ---------------*
.subckt PWR_CHNEL_1 A1 A2 VPB VPWR Y2 W1=4 L1=1 W2=4 L2=1
XM1_BIAS1_f1 Y1 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w="W1" l="L1"
XM1_BIAS2_f1 Y2 A2 Y1 VPB sky130_fd_pr__pfet_01v8_hvt	 w="W2" l="L2"
.ends

.subckt PWR_CHNEL_2 A1 A2 VPB VPWR Y2 W1=4 L1=1 W2=4 L2=1
XM1_BIAS1_f1 Y1 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w="W1" l="L1"
XM1_BIAS1_f2 VPWR A1 Y1 VPB sky130_fd_pr__pfet_01v8_hvt w="W1" l="L1"
XM1_BIAS2_f1 Y2 A2 Y1 VPB sky130_fd_pr__pfet_01v8_hvt  w="W2" l="L2"
XM1_BIAS2_f2 Y1 A2 Y2 VPB sky130_fd_pr__pfet_01v8_hvt  w="W2" l="L2
.ends

.subckt I_LOCK KEY ADD_PWR VGND VNB VPB VPWR I_SUP 
+ Wp_lk=4 Lp_lk=1 Wn_lk=2 Ln_lk=1 Wp_op=4 Lp_op=1 Wn_op=2 Ln_op=1 Rl=100
X_inv_1 KEY VGND VNB VPB VPWR KEY_INV sky130_fd_sc_hd__inv_2
** Lock 
XMp_lk_f1 ADD_PWR KEY rLOAD VPB sky130_fd_pr__pfet_01v8 		w="Wp_lk" l="Lp_lk"
XMp_lk_f2 rLOAD KEY ADD_PWR VPB sky130_fd_pr__pfet_01v8 		w="Wp_lk" l="Lp_lk"
XMn_lk_f1 ADD_PWR KEY_INV rLOAD VNB sky130_fd_pr__nfet_01v8 w="Wn_lk" l="Ln_lk"
XMn_lk_f2 rLOAD KEY_INV ADD_PWR VNB sky130_fd_pr__nfet_01v8 w="Wn_lk" l="Ln_lk"
R_dsch rLOAD GND R={Rl}
** Open
XMp_op_f1 ADD_PWR KEY_INV I_SUP VPB sky130_fd_pr__pfet_01v8 w="Wp_op" l="Lp_op"
XMp_op_f2 I_SUP KEY_INV ADD_PWR VPB sky130_fd_pr__pfet_01v8 w="Wp_op" l="Lp_op"
XMn_op_f1 ADD_PWR KEY I_SUP VNB sky130_fd_pr__nfet_01v8 		w="Wn_op" l="Ln_op"
XMn_op_f2 I_SUP KEY ADD_PWR VNB sky130_fd_pr__nfet_01v8 		w="Wn_op" l="Ln_op"
.ends

.subckt I_DAC KEY V_BIAS1 V_BIAS2 V_BIAS3 V_BIAS4 VGND VNB VPB VPWR I_SUP 	$INTERNAL 1-BIT DAC SUB CIRCUIT
+ W_br1=4 L_br1=1 W_br2=4 L_br2=1
+ Wp_lk=4 Lp_lk=1 Wn_lk=2 Ln_lk=1 Rl=100
X_BRAN_1 V_BIAS1 V_BIAS2 VPB VPWR I_SUP	$ Branch_1 Transistors Power Supply (maintain)
+ PWR_CHNEL_1 W1="W_br1" L1="L_br1" W2="W_br1" L2="L_br1"
X_BRAN_2 V_BIAS3 V_BIAS4 VPB VPWR ADD_PWR    $ Branch_2 Transistors Power Supply (addition)
+ PWR_CHNEL_2 W1="W_br2" L1="L_br2" W2="W_br2" L2="L_br2"
X_LOCK KEY ADD_PWR VGND VNB VPB VPWR I_SUP I_LOCK		$ Digital Control Block
+ Wp_lk="Wp_lk" Lp_lk="Lp_lk" Wn_lk="Wn_lk" Ln_lk="Ln_lk"
+ Wp_op="Wp_lk" Lp_op="Lp_lk" Wn_op="Wn_lk" Ln_op="Ln_lk" Rl="Rl"
.ends

.subckt FREQ_DIV2 CLK VGND VNB VPB VPWR CLK_DIV2_buf   $ FREQUENCY DIVIDER
X_buffer1 CLK VGND VNB VPB VPWR CLK_BUF sky130_fd_sc_ms__clkbuf_2
X_STAGE1 CLK_BUF D1 VGND VNB VPB VPWR CLK_DIV2 Q1N sky130_fd_sc_ms__dfxbp_1
X_dly1 Q1N VGND VNB VPB VPWR DL1 sky130_fd_sc_ms__dlygate4sd3_1
X_dly2 DL1 VGND VNB VPB VPWR DL2 sky130_fd_sc_ms__dlygate4sd3_1
X_dly3 DL2 VGND VNB VPB VPWR DL3 sky130_fd_sc_ms__dlygate4sd3_1
X_dly4 DL3 VGND VNB VPB VPWR DL4 sky130_fd_sc_ms__dlygate4sd3_1
X_dly5 DL4 VGND VNB VPB VPWR Dl5 sky130_fd_sc_ms__dlygate4sd3_1
X_dly6 DL5 VGND VNB VPB VPWR D1 sky130_fd_sc_ms__dlygate4sd3_1
X_buffer2 CLK_DIV2 VGND VNB VPB VPWR CLK_DIV2_buf sky130_fd_sc_ms__clkbuf_1
.ends

.subckt CAP_ARR NDp[0] NDp[1] NDp[2] NDp[3] NDp[4] NDn[0] NDn[1] NDn[2] NDn[3] NDn[4] Cap="Cap"
C1p NDp[0] gnd C=Cap 		$ CAPACITOR ARRAY
C2p NDp[1] gnd C=Cap
C3p NDp[2] gnd C=Cap
C4p NDp[3] gnd C=Cap
C5p NDp[4] gnd C=Cap
C1n NDn[0] gnd C=Cap
C2n NDn[1] gnd C=Cap
C3n NDn[2] gnd C=Cap
C4n NDn[3] gnd C=Cap
C5n NDn[4] gnd C=Cap
.ends

.subckt VCO_STARTUP ENB VGND VNB VPB VPWR START_PWL 
* STARTUP OSCILLATION
Xconb_1 VGND VNB VPB VPWR hi_logic lo_logic sky130_fd_sc_hd__conb_1
Xeinvp_1 hi_logic ENB VGND VNB VPB VPWR p[0] sky130_fd_sc_hd__einvp_1
.ends

*****----------*****----------*****----------*****----------*****----------*****
*
*_____________DCO design process__________________*
* RING_OSC-1
Xr1 p[0] p[1] p[2] p[3] p[4] p_n[0] p_n[1] p_n[2] p_n[3] p_n[4]
+ gnd gnd I_SUP I_SUP ring_osc_s1
+ Wp12=Wp12 Wn12=Wn12 L12=L12
+ Wp34=Wp34 Wn34=Wn34 L34=L34

* X_STARTUP ENB GND GND VDD VDD str VCO_STARTUP

*X_CapArr p[0] p[1] p[2] p[3] p[4] p_n[0] p_n[1] p_n[2] p_n[3] p_n[4] CAP_ARR Cap=C_insert $ CAPACITOR ARRAY

X_DAC D_1 Vbs1 Vbs2 Vbs3 Vbs4 gnd gnd VCA VCA load I_DAC 	$ INTERNAL 1-BIT DAC
+ W_br1=W_br1  L_br1=L_br1  W_br2=W_br2  L_br2=L_br2
+ Wp_lk=Wp_lk  Lp_lk=Lp_lk  Wn_lk=Wn_lk  Ln_lk=Ln_lk Rl=50000

X_CLK_DIV2 p[0] gnd gnd VCD VCD CLK_DIV2 FREQ_DIV2 	$ FREQUENCY DIVIDER

*********************************************
** Debug zone **

R_debug load I_SUP R=0.01
* VOLTAGE REFERENCE
Vsup V_sup gnd DC=1.8
V_a VCA gnd	DC=1.8
V_d VCD gnd	DC=1.8
V2 Vbs1 gnd DC=0.3
V3 Vbs2 gnd DC=0.3
V4 Vbs3 gnd DC=0
V5 Vbs4 gnd DC=0
V6 ENB  gnd DC=0 PULSE( 0 1.8 0 20n 20n 200n 1 )
V7 D_1  gnd DC=1.8 $PULSE( 0 1.8 0 0.2n 0.2n 2u 5u )
V8 CLK  gnd DC=0 PULSE( 0 1.8 0 2n 2n 18n 40n ) 

***-------parameters--------***
.param W_br1=1
.param L_br1=0.5
.param W_br2=2.4
.param L_br2=0.5
.param Wp_lk=4
.param Lp_lk=0.5
.param Wn_lk=2
.param Ln_lk=0.5
 
.param Wp12=5
.param Wn12=2
.param L12=2
.param Wp34=2.5
.param Wn34=1
.param L34=2
*.param C_insert= 15f

* CONTROL TESTBENCH
.control 
set test_mode = 2
set num_threads = 8
** mode = 0:operation testing * 1:frequency extract * 2:power consumption *3:generate data 
*
if ($test_mode = 2) 
	save @R_debug[i] "p[0]" load I_SUP @V_a[i] VCA CLK_DIV2 CLK_BUF D1 D2
	TRAN 1n 16u
	MEAS TRAN I_osc AVG @R_debug[i] FROM=4u TO=10u
	MEAS TRAN I_dco1 AVG @V_a[i] FROM=4u TO=10u
	MEAS TRAN V_dco AVG VCA FROM=4u TO=10u
	MEAS TRAN prd TRIG CLK_DIV2 VAL=0.8 RISE=10 TARG CLK_DIV2 VAL=0.8 RISE=30
	let Power_f = I_dco1*V_dco	
	let freq = 20/prd
	plot "p[0]" clk_div2
*	plot @V1[i]
	print freq I_dco1 I_osc Power_f
end 

if ($test_mode = 0)
	TRAN 1n 6u
	plot "p[0]" CLK_DIV4
	MEAS TRAN prd TRIG p[0] VAL=0.8 RISE=5 TARG p[0] VAL=0.8 RISE=25
	MEAS TRAN prd1 TRIG CLK_DIV4 VAL=0.8 RISE=5 TARG CLK_DIV4 VAL=0.8 RISE=10
	MEAS TRAN I_dco AVG @V1[i] FROM=2u TO=5u
	let freq = 20/prd
	let freq_div4 = 5/prd1
	echo "frequency: " 
	print freq freq_div4 I_dco
end 

if ($test_mode = 1)
	let Vlow = 1.19			$ set lower bound for sweeping 
	let Vlimit = 1.8		$ set upper bound for sweeping
	let Vsweep = 0.2		$ set step size for sweeping
	let NoPoints=(Vlimit-Vlow)/Vsweep+2		$ set number of points for sweeping
	let freq =unitvec(NoPoints)
	let freq_div2 =unitvec(NoPoints)
	let Vin  =unitvec(NoPoints)
	let Vosc =unitvec(NoPoints)
	let Iosc =unitvec(NoPoints)
	let Power=unitvec(NoPoints)
	let Vin[0]=Vlimit
	let ix=0
	save V_sup @Vsup[i] "p[0]" Wp12 Wn12 Wp34 Wn34 L12 L34 enb CLK_DIV4 clk_div2
	while Vin[ix] > Vlow
		alter Vsup DC=Vin[ix]
		if Vin[ix] < 1.5
			TRAN 0.5n 12u
		else
			TRAN 0.5n 5u
		end
		MEAS TRAN prd TRIG p[0] VAL=0.8 RISE=5 TARG p[0] VAL=0.8 RISE =15
		MEAS TRAN prd1 TRIG CLK_DIV2 VAL=0.8 RISE=5 TARG CLK_DIV2 VAL=0.8 RISE =15
		MEAS TRAN I_vco AVG @Vsup[i] FROM=1u TO=2u
		MEAS TRAN V_vco AVG V_sup FROM=1u TO=2u
		let freq[ix] = 10/prd
		let freq_div2[ix] = 10/prd1
		let Power[ix]=I_vco*V_vco
		let Iosc[ix]=I_vco
		let ix = ix+1
		Let Vin[ix] = Vin[ix-1]-Vsweep
	end	
	print Vin freq freq_div2 power Iosc
	plot "p[0]" CLK_DIV2
end

.endc
