magic
tech sky130A
timestamp 1723779942
<< nwell >>
rect 270 640 350 660
rect 900 640 980 660
rect 230 620 390 640
rect 870 630 1030 640
rect 180 510 250 540
rect 260 520 380 620
rect 260 480 370 520
rect 830 500 860 530
rect 260 470 360 480
rect 180 430 250 470
rect 270 400 360 470
rect 900 420 990 630
rect 270 290 350 400
rect 560 380 590 410
rect 900 290 980 420
rect 1360 380 1390 410
<< pwell >>
rect 270 170 350 250
rect 250 0 360 170
rect 900 0 980 250
rect 1100 150 1140 200
rect 1360 120 1390 150
<< nmos >>
rect 1100 150 1140 200
<< ndiffc >>
rect 1360 120 1390 150
<< pdiffc >>
rect 830 500 860 530
rect 200 440 230 470
rect 560 380 590 410
rect 1360 380 1390 410
<< psubdiff >>
rect 290 60 340 80
rect 290 30 300 60
rect 330 30 340 60
rect 290 10 340 30
rect 920 60 970 80
rect 920 30 930 60
rect 960 30 970 60
rect 920 10 970 30
<< nsubdiff >>
rect 290 600 340 620
rect 290 570 300 600
rect 330 570 340 600
rect 290 550 340 570
rect 920 590 970 610
rect 920 560 930 590
rect 960 560 970 590
rect 920 540 970 560
rect 290 390 340 410
rect 290 360 300 390
rect 330 360 340 390
rect 290 340 340 360
<< psubdiffcont >>
rect 300 30 330 60
rect 930 30 960 60
<< nsubdiffcont >>
rect 300 570 330 600
rect 930 560 960 590
rect 300 360 330 390
<< poly >>
rect 10 280 90 290
rect 1170 280 1240 290
rect 30 260 50 280
rect 70 260 90 280
rect 1190 260 1210 280
rect 1230 260 1240 280
rect 10 250 90 260
rect 1170 250 1240 260
<< polycont >>
rect -70 260 -50 280
rect -30 260 -10 280
rect 10 260 30 280
rect 50 260 70 280
rect 90 260 110 280
rect 130 260 150 280
rect 460 260 480 280
rect 500 260 520 280
rect 730 260 750 280
rect 770 260 790 280
rect 1090 260 1110 280
rect 1130 260 1150 280
rect 1170 260 1190 280
rect 1210 260 1230 280
rect 1250 260 1270 280
rect 1290 260 1310 280
<< locali >>
rect 290 600 340 620
rect 290 570 300 600
rect 330 570 340 600
rect 920 590 970 610
rect 290 390 340 570
rect 920 560 930 590
rect 960 560 970 590
rect 920 540 970 560
rect 290 360 300 390
rect 330 360 340 390
rect 290 340 340 360
rect -90 280 180 290
rect -90 260 -70 280
rect -50 260 -30 280
rect -10 260 10 280
rect 30 260 50 280
rect 70 260 90 280
rect 110 260 130 280
rect 150 260 180 280
rect -90 250 180 260
rect 210 230 250 310
rect 440 280 540 290
rect 440 260 460 280
rect 480 260 500 280
rect 520 260 540 280
rect 440 250 540 260
rect 570 230 610 310
rect 710 280 810 290
rect 710 260 730 280
rect 750 260 770 280
rect 790 260 810 280
rect 710 250 810 260
rect 840 230 880 310
rect 1070 280 1340 290
rect 1070 260 1090 280
rect 1110 260 1130 280
rect 1150 260 1170 280
rect 1190 260 1210 280
rect 1230 260 1250 280
rect 1270 260 1290 280
rect 1310 260 1340 280
rect 1070 250 1340 260
rect 1370 230 1410 310
rect 290 60 340 80
rect 290 30 300 60
rect 330 30 340 60
rect 290 10 340 30
rect 920 60 970 80
rect 920 30 930 60
rect 960 30 970 60
rect 920 10 970 30
<< viali >>
rect -140 560 -110 590
rect 300 570 330 600
rect 200 500 230 530
rect 200 440 230 470
rect 390 560 420 590
rect 660 560 690 590
rect 930 560 960 590
rect 1020 560 1050 590
rect 830 500 860 530
rect 830 440 860 470
rect 300 360 330 390
rect 560 380 590 410
rect 1360 380 1390 410
rect 200 330 230 360
rect 560 330 590 360
rect 1360 330 1390 360
rect -70 260 -50 280
rect -30 260 -10 280
rect 10 260 30 280
rect 50 260 70 280
rect 90 260 110 280
rect 130 260 150 280
rect 460 260 480 280
rect 500 260 520 280
rect 730 260 750 280
rect 770 260 790 280
rect 1090 260 1110 280
rect 1130 260 1150 280
rect 1170 260 1190 280
rect 1210 260 1230 280
rect 1250 260 1270 280
rect 1290 260 1310 280
rect 200 180 230 210
rect 560 180 590 210
rect 1360 180 1390 210
rect 1360 120 1390 150
rect 300 30 330 60
rect 930 30 960 60
<< metal1 >>
rect -160 590 -90 700
rect -160 560 -140 590
rect -110 560 -90 590
rect -160 545 -90 560
rect 290 600 340 620
rect 290 570 300 600
rect 330 570 340 600
rect 290 550 340 570
rect 370 590 440 700
rect 370 560 390 590
rect 420 560 440 590
rect 370 545 440 560
rect 640 590 710 700
rect 640 560 660 590
rect 690 560 710 590
rect 640 545 710 560
rect 920 590 970 610
rect 920 560 930 590
rect 960 560 970 590
rect 920 540 970 560
rect 1000 590 1070 700
rect 1000 560 1020 590
rect 1050 560 1070 590
rect 1000 545 1070 560
rect 180 530 250 540
rect -180 470 -20 510
rect -60 290 -20 470
rect 180 500 200 530
rect 230 510 250 530
rect 810 530 880 540
rect 810 510 830 530
rect 230 500 830 510
rect 860 510 880 530
rect 860 500 1430 510
rect 180 470 1430 500
rect 180 440 200 470
rect 230 440 250 470
rect 180 430 250 440
rect 810 440 830 470
rect 860 440 880 470
rect 810 430 880 440
rect 540 410 610 420
rect 290 390 340 410
rect 180 360 250 370
rect 180 330 200 360
rect 230 330 250 360
rect 290 360 300 390
rect 330 360 340 390
rect 290 340 340 360
rect 540 380 560 410
rect 590 380 610 410
rect 540 370 610 380
rect 1340 410 1410 420
rect 1340 380 1360 410
rect 1390 380 1410 410
rect 1340 370 1410 380
rect 540 360 1410 370
rect 180 310 250 330
rect 540 330 560 360
rect 590 330 1360 360
rect 1390 330 1410 360
rect 540 310 610 330
rect 210 290 250 310
rect 570 290 610 310
rect 740 290 780 330
rect 1340 310 1410 330
rect -90 280 180 290
rect -90 260 -70 280
rect -50 260 -30 280
rect -10 260 10 280
rect 30 260 50 280
rect 70 260 90 280
rect 110 260 130 280
rect 150 260 180 280
rect -90 250 180 260
rect 210 280 540 290
rect 210 260 460 280
rect 480 260 500 280
rect 520 260 540 280
rect 210 250 540 260
rect 570 280 810 290
rect 570 260 730 280
rect 750 260 770 280
rect 790 260 810 280
rect 570 250 810 260
rect 1070 280 1340 290
rect 1070 260 1090 280
rect 1110 260 1130 280
rect 1150 260 1170 280
rect 1190 260 1210 280
rect 1230 260 1250 280
rect 1270 260 1290 280
rect 1310 260 1340 280
rect 1070 250 1340 260
rect 210 230 250 250
rect 570 230 610 250
rect 180 210 250 230
rect 180 180 200 210
rect 230 180 250 210
rect 180 170 250 180
rect 540 210 610 230
rect 540 180 560 210
rect 590 180 610 210
rect 540 170 610 180
rect 1100 150 1140 250
rect -180 110 1140 150
rect 1340 210 1410 230
rect 1340 180 1360 210
rect 1390 180 1410 210
rect 1340 150 1410 180
rect 1340 120 1360 150
rect 1390 120 1430 150
rect 1340 110 1430 120
rect 290 60 340 80
rect 290 30 300 60
rect 330 30 340 60
rect 290 10 340 30
rect 920 60 970 80
rect 920 30 930 60
rect 960 30 970 60
rect 920 10 970 30
use inv_d  inv_d_0
timestamp 1723626483
transform 1 0 80 0 1 310
box -90 -310 190 350
use inv_d  inv_d_1
timestamp 1723626483
transform 1 0 440 0 1 310
box -90 -310 190 350
use inv_d  inv_d_2
timestamp 1723626483
transform 1 0 710 0 1 310
box -90 -310 190 350
use inv_d  inv_d_3
timestamp 1723626483
transform 1 0 1070 0 1 310
box -90 -310 190 350
use inv_d  inv_d_4
timestamp 1723626483
transform 1 0 -90 0 1 310
box -90 -310 190 350
use inv_d  inv_d_5
timestamp 1723626483
transform 1 0 1240 0 1 310
box -90 -310 190 350
<< labels >>
rlabel metal1 -180 490 -180 490 7 inp
port 1 w
rlabel metal1 -180 130 -180 130 7 inn
port 2 w
rlabel metal1 1430 490 1430 490 3 outp
port 3 e
rlabel metal1 1430 130 1430 130 3 outn
port 4 e
<< end >>
