magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 523 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 129 247 177
rect 193 95 203 129
rect 237 95 247 129
rect 193 47 247 95
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 129 415 177
rect 361 95 371 129
rect 405 95 415 129
rect 361 47 415 95
rect 445 161 497 177
rect 445 127 455 161
rect 489 127 497 161
rect 445 93 497 127
rect 445 59 455 93
rect 489 59 497 93
rect 445 47 497 59
<< pdiff >>
rect 27 479 79 497
rect 27 445 35 479
rect 69 445 79 479
rect 27 411 79 445
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 463 247 497
rect 193 429 203 463
rect 237 429 247 463
rect 193 368 247 429
rect 193 334 203 368
rect 237 334 247 368
rect 193 297 247 334
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 297 331 383
rect 361 463 415 497
rect 361 429 371 463
rect 405 429 415 463
rect 361 368 415 429
rect 361 334 371 368
rect 405 334 415 368
rect 361 297 415 334
rect 445 485 497 497
rect 445 451 455 485
rect 489 451 497 485
rect 445 417 497 451
rect 445 383 455 417
rect 489 383 497 417
rect 445 349 497 383
rect 445 315 455 349
rect 489 315 497 349
rect 445 297 497 315
<< ndiffc >>
rect 35 95 69 129
rect 119 63 153 97
rect 203 95 237 129
rect 287 63 321 97
rect 371 95 405 129
rect 455 127 489 161
rect 455 59 489 93
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 119 451 153 485
rect 119 383 153 417
rect 203 429 237 463
rect 203 334 237 368
rect 287 451 321 485
rect 287 383 321 417
rect 371 429 405 463
rect 371 334 405 368
rect 455 451 489 485
rect 455 383 489 417
rect 455 315 489 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 79 261 109 297
rect 28 249 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 415 259 445 297
rect 28 215 44 249
rect 78 215 109 249
rect 28 203 109 215
rect 162 249 445 259
rect 162 215 178 249
rect 212 215 445 249
rect 162 205 445 215
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 177 445 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
<< polycont >>
rect 44 215 78 249
rect 178 215 212 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 485 167 527
rect 153 451 167 485
rect 119 417 167 451
rect 153 383 167 417
rect 119 367 167 383
rect 203 463 237 493
rect 203 368 237 429
rect 19 309 35 343
rect 69 331 85 343
rect 271 485 337 527
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 271 367 337 383
rect 371 463 405 493
rect 371 368 405 429
rect 69 309 162 331
rect 19 297 162 309
rect 18 249 94 263
rect 18 215 44 249
rect 78 215 94 249
rect 128 249 162 297
rect 203 323 237 334
rect 371 323 405 334
rect 203 289 405 323
rect 439 485 505 527
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 439 349 505 383
rect 439 315 455 349
rect 489 315 505 349
rect 439 297 505 315
rect 128 215 178 249
rect 212 215 228 249
rect 128 181 162 215
rect 306 181 405 289
rect 35 147 162 181
rect 203 147 405 181
rect 35 129 69 147
rect 203 129 237 147
rect 35 51 69 95
rect 105 97 153 113
rect 105 63 119 97
rect 105 17 153 63
rect 371 129 405 147
rect 203 51 237 95
rect 271 97 337 113
rect 271 63 287 97
rect 321 63 337 97
rect 271 17 337 63
rect 371 51 405 95
rect 439 161 505 177
rect 439 127 455 161
rect 489 127 505 161
rect 439 93 505 127
rect 439 59 455 93
rect 489 59 505 93
rect 439 17 505 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 X
port 4 nsew
flabel locali s 306 289 340 323 0 FreeSans 200 0 0 0 X
port 4 nsew
flabel locali s 306 153 340 187 0 FreeSans 200 0 0 0 X
port 4 nsew
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 5 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew
rlabel comment s 0 0 0 0 4 buf_4
<< properties >>
string FIXED_BBOX 0 0 552 544
string path 0.000 2.720 2.760 2.720 
<< end >>
