magic
tech sky130A
magscale 1 2
timestamp 1727163546
<< nwell >>
rect 3080 3500 3256 3820
rect 7210 900 7340 1220
<< pwell >>
rect 3156 3258 3290 3394
rect 7170 660 7340 840
<< psubdiff >>
rect 3178 3342 3240 3376
rect 3178 3308 3194 3342
rect 3230 3308 3240 3342
rect 3178 3276 3240 3308
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7230 700 7290 730
<< nsubdiff >>
rect 3160 3662 3220 3696
rect 3160 3628 3174 3662
rect 3208 3628 3220 3662
rect 3160 3596 3220 3628
rect 7230 1020 7290 1050
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
<< psubdiffcont >>
rect 3194 3308 3230 3342
rect 7240 730 7280 770
<< nsubdiffcont >>
rect 3174 3628 3208 3662
rect 7240 980 7280 1020
<< locali >>
rect 3160 3670 3220 3696
rect 3730 3670 4190 3730
rect 3160 3630 3170 3670
rect 3210 3630 3220 3670
rect 3160 3628 3174 3630
rect 3208 3628 3220 3630
rect 3160 3596 3220 3628
rect 3690 3490 3760 3500
rect 3690 3450 3700 3490
rect 3740 3450 3760 3490
rect 3690 3440 3760 3450
rect 3170 3342 3240 3380
rect 3170 3308 3194 3342
rect 3230 3308 3240 3342
rect 3170 3170 3240 3308
rect 3290 3170 3360 3230
rect 3170 3100 3360 3170
rect 3170 2730 3270 3100
rect 4130 3040 4190 3670
rect 4400 3440 5390 3460
rect 4400 3400 5330 3440
rect 5370 3400 5390 3440
rect 4400 3380 5390 3400
rect 4120 3020 4200 3040
rect 4120 2980 4140 3020
rect 4180 2980 4200 3020
rect 4120 2960 4200 2980
rect 4400 2730 4480 3380
rect 3170 2650 4480 2730
rect 3170 1020 3270 2650
rect 3170 970 3190 1020
rect 3240 970 3270 1020
rect 3170 940 3270 970
rect 5980 1540 6080 1560
rect 5980 1500 6010 1540
rect 6050 1500 6080 1540
rect 2160 600 2340 680
rect 5980 -270 6080 1500
rect 7950 1360 8460 1390
rect 7950 1320 7980 1360
rect 8020 1320 8060 1360
rect 8100 1320 8140 1360
rect 8180 1320 8220 1360
rect 8260 1320 8300 1360
rect 8340 1320 8380 1360
rect 8420 1320 8460 1360
rect 7950 1290 8460 1320
rect 7230 1020 7290 1050
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7090 490 7170 630
rect 7230 490 7290 730
rect 7090 430 7290 490
rect 7950 480 8050 1290
rect 8360 630 8460 1290
rect 7090 250 7170 430
rect 7090 150 7620 250
rect 7090 110 7190 150
rect 8410 110 8440 120
rect 7090 30 8440 110
rect 7090 -2090 7190 30
rect 7090 -2190 7620 -2090
rect 7090 -2230 7190 -2190
rect 8410 -2230 8450 -2220
rect 7090 -2300 8450 -2230
rect 2750 -4080 2950 -3120
rect 7090 -4080 7190 -2300
rect 2750 -4280 7420 -4080
<< viali >>
rect 2600 5860 2640 5900
rect 3180 5860 3220 5900
rect 3760 5860 3800 5900
rect 4620 5860 4660 5900
rect 5480 5860 5520 5900
rect 6060 5860 6100 5900
rect 6640 5860 6680 5900
rect 7500 5860 7540 5900
rect 8360 5860 8400 5900
rect 8940 5860 8980 5900
rect 9520 5860 9560 5900
rect 2600 4200 2640 4240
rect 3180 4200 3220 4240
rect 3760 4200 3800 4240
rect 4620 4200 4660 4240
rect 5480 4200 5520 4240
rect 6060 4200 6100 4240
rect 6640 4200 6680 4240
rect 7500 4200 7540 4240
rect 8360 4200 8400 4240
rect 8940 4200 8980 4240
rect 3170 3662 3210 3670
rect 3170 3630 3174 3662
rect 3174 3630 3208 3662
rect 3208 3630 3210 3662
rect 3330 3460 3370 3500
rect 3700 3450 3740 3490
rect 3194 3308 3230 3342
rect 5330 3400 5370 3440
rect 5910 3400 5950 3440
rect 6490 3400 6530 3440
rect 7350 3400 7390 3440
rect 8210 3400 8250 3440
rect 8790 3400 8830 3440
rect 9370 3400 9410 3440
rect 4140 2980 4180 3020
rect 5330 1740 5370 1780
rect 5910 1740 5950 1780
rect 6490 1740 6530 1780
rect 7350 1740 7390 1780
rect 8210 1740 8250 1780
rect 8790 1740 8830 1780
rect 9370 1740 9410 1780
rect 10230 1740 10270 1780
rect 3190 970 3240 1020
rect 6010 1500 6050 1540
rect 7980 1320 8020 1360
rect 8060 1320 8100 1360
rect 8140 1320 8180 1360
rect 8220 1320 8260 1360
rect 8300 1320 8340 1360
rect 8380 1320 8420 1360
rect 7028 1050 7062 1084
rect 7028 974 7062 1008
rect 7240 980 7280 1020
rect 6846 854 6880 888
rect 7240 730 7280 770
<< metal1 >>
rect 4520 5340 4740 5420
rect 3160 3820 3300 3830
rect 3160 3760 3170 3820
rect 3230 3760 3300 3820
rect 3160 3740 3300 3760
rect 3920 3810 4010 3830
rect 3920 3750 3940 3810
rect 4000 3750 4010 3810
rect 3160 3670 3220 3740
rect 3160 3630 3170 3670
rect 3210 3630 3220 3670
rect 3160 3596 3220 3630
rect 3300 3500 3400 3540
rect 3920 3500 4010 3750
rect 3300 3490 3330 3500
rect 2890 3460 3330 3490
rect 3370 3460 3400 3500
rect 2890 3430 3400 3460
rect 3680 3490 4010 3500
rect 3680 3450 3700 3490
rect 3740 3450 4010 3490
rect 3680 3430 4010 3450
rect 3178 3342 3240 3376
rect 3178 3308 3194 3342
rect 3230 3308 3240 3342
rect 3178 3276 3240 3308
rect 4220 1240 4300 2280
rect 7180 1380 7290 1390
rect 7180 1320 7210 1380
rect 7270 1320 7290 1380
rect 4220 1160 6490 1240
rect 7180 1230 7290 1320
rect 7950 1370 8460 1390
rect 7950 1310 7970 1370
rect 8030 1360 8130 1370
rect 8190 1360 8290 1370
rect 8350 1360 8460 1370
rect 8030 1320 8060 1360
rect 8100 1320 8130 1360
rect 8190 1320 8220 1360
rect 8260 1320 8290 1360
rect 8350 1320 8380 1360
rect 8420 1320 8460 1360
rect 8030 1310 8130 1320
rect 8190 1310 8290 1320
rect 8350 1310 8460 1320
rect 7950 1290 8460 1310
rect 3170 1020 6270 1040
rect 3170 970 3190 1020
rect 3240 970 6270 1020
rect 2540 870 2640 960
rect 3170 940 6270 970
rect 2540 770 5590 870
rect 2540 480 2640 770
rect 3960 480 4060 590
rect 3750 380 4390 480
rect 5490 470 5590 770
rect 6170 250 6270 940
rect 6410 910 6490 1160
rect 7160 1140 7290 1230
rect 7020 1084 7070 1100
rect 7020 1050 7028 1084
rect 7062 1050 7070 1084
rect 7020 1008 7070 1050
rect 7020 974 7028 1008
rect 7062 974 7070 1008
rect 6410 908 6830 910
rect 6410 888 6896 908
rect 6410 854 6846 888
rect 6880 854 6896 888
rect 7020 900 7070 974
rect 7230 1020 7290 1140
rect 7230 980 7240 1020
rect 7280 980 7290 1020
rect 7230 950 7290 980
rect 7350 900 8270 930
rect 7020 860 8270 900
rect 7037 858 8270 860
rect 6410 836 6896 854
rect 6410 830 6830 836
rect 7350 830 8270 858
rect 7230 770 7290 800
rect 7230 730 7240 770
rect 7280 730 7290 770
rect 7230 700 7290 730
rect 8170 350 8270 830
rect 6170 150 7540 250
rect 11080 -70 11180 -50
rect 11080 -130 11100 -70
rect 11160 -130 11180 -70
rect 11080 -150 11180 -130
rect 11840 -70 11940 -50
rect 11840 -130 11860 -70
rect 11920 -130 11940 -70
rect 1240 -1540 1320 -1340
rect 1540 -1360 1640 -1340
rect 1540 -1420 1560 -1360
rect 1620 -1420 1640 -1360
rect 1540 -1480 1640 -1420
rect 11840 -1430 11940 -130
rect 8140 -1530 11940 -1430
rect 6530 -1780 7730 -1760
rect 6530 -1840 6550 -1780
rect 6610 -1840 7730 -1780
rect 6530 -1860 7730 -1840
rect 8040 -1860 8050 -1760
rect 8140 -1960 8240 -1530
rect 11080 -2410 11180 -2390
rect 11080 -2470 11100 -2410
rect 11160 -2470 11180 -2410
rect 7680 -2580 7930 -2490
rect 11080 -2500 11180 -2470
<< via1 >>
rect 3170 3760 3230 3820
rect 3940 3750 4000 3810
rect 7210 1320 7270 1380
rect 7970 1360 8030 1370
rect 8130 1360 8190 1370
rect 8290 1360 8350 1370
rect 7970 1320 7980 1360
rect 7980 1320 8020 1360
rect 8020 1320 8030 1360
rect 8130 1320 8140 1360
rect 8140 1320 8180 1360
rect 8180 1320 8190 1360
rect 8290 1320 8300 1360
rect 8300 1320 8340 1360
rect 8340 1320 8350 1360
rect 7970 1310 8030 1320
rect 8130 1310 8190 1320
rect 8290 1310 8350 1320
rect 11100 -130 11160 -70
rect 11860 -130 11920 -70
rect 1560 -1420 1620 -1360
rect 6550 -1840 6610 -1780
rect 11100 -2470 11160 -2410
<< metal2 >>
rect -720 3830 -530 6080
rect -720 3820 4010 3830
rect -720 3760 3170 3820
rect 3230 3810 4010 3820
rect 3230 3760 3940 3810
rect -720 3750 3940 3760
rect 4000 3750 4010 3810
rect -720 3740 4010 3750
rect -720 1390 -530 3740
rect -720 1380 8460 1390
rect -720 1320 7210 1380
rect 7270 1370 8460 1380
rect 7270 1320 7970 1370
rect -720 1310 7970 1320
rect 8030 1310 8130 1370
rect 8190 1310 8290 1370
rect 8350 1310 8460 1370
rect -720 1300 8460 1310
rect -720 145 -530 1300
rect 1540 -1360 1640 1300
rect 1540 -1420 1560 -1360
rect 1620 -1420 1640 -1360
rect 1540 -1440 1640 -1420
rect 6530 -1780 6630 1300
rect 7950 1290 8460 1300
rect 11080 -70 11940 -50
rect 11080 -130 11100 -70
rect 11160 -130 11860 -70
rect 11920 -130 11940 -70
rect 11080 -150 11940 -130
rect 6530 -1840 6550 -1780
rect 6610 -1840 6630 -1780
rect 6530 -1860 6630 -1840
rect 11080 -2410 11890 -2390
rect 11080 -2470 11100 -2410
rect 11160 -2470 11890 -2410
rect 11080 -2490 11890 -2470
use dco_freq  dco_freq_0
timestamp 1726743291
transform 1 0 8320 0 1 50
box -880 -1250 3330 640
use dco_freq  dco_freq_1
timestamp 1726743291
transform 1 0 8320 0 1 -2290
box -880 -1250 3330 640
use dco_idac  dco_idac_0
timestamp 1727082698
transform 1 0 2860 0 1 -60
box -1860 -3160 3220 740
use dco_ring_osc  dco_ring_osc_0
timestamp 1726107115
transform 1 0 1680 0 1 4000
box -500 -2520 9440 2160
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 6808 0 1 638
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 3288 0 1 3238
box -38 -48 498 592
<< labels >>
rlabel locali 6040 1560 6040 1560 1 Isup
rlabel metal1 4010 590 4010 590 1 Vbs_34
port 6 n
rlabel metal1 2590 960 2590 960 1 Vbs_12
port 5 n
rlabel metal2 11900 -50 11900 -50 1 ro_div2
rlabel metal2 11820 -2390 11820 -2390 1 pha_DCO
port 7 n
rlabel metal1 7560 930 7560 930 1 pha_ro
rlabel metal1 4340 1240 4340 1240 1 p_osc
rlabel metal2 -620 6080 -620 6080 1 VCCD
port 1 n
rlabel metal1 2930 3490 2930 3490 1 ENB
port 4 n
rlabel locali 2190 680 2190 680 1 VCCA
port 2 n
rlabel metal1 1290 -1340 1290 -1340 1 Dctrl
port 3 n
rlabel locali 4910 -4080 4910 -4080 1 GND
port 8 n
<< end >>
