magic
tech sky130A
magscale 1 2
timestamp 1724225882
<< pwell >>
rect 3990 1550 4520 1810
<< locali >>
rect 3410 2510 3510 3060
rect 3740 2000 3820 2030
rect 3740 1960 3760 2000
rect 3800 1960 3820 2000
rect 3740 1700 3820 1960
rect 3740 1620 4050 1700
rect 3990 1540 4090 1560
rect 3990 1500 4020 1540
rect 4060 1500 4090 1540
rect 3990 1470 4090 1500
<< viali >>
rect 3760 1960 3800 2000
rect 4020 1500 4060 1540
rect 4410 1500 4450 1540
rect 4410 1420 4450 1460
<< metal1 >>
rect 2170 3210 2270 3560
rect 850 3130 950 3210
rect 2100 3130 2270 3210
rect 2170 2590 2270 3130
rect 2170 2510 2310 2590
rect 3390 1540 4090 1570
rect 3390 1500 4020 1540
rect 4060 1500 4090 1540
rect 3390 1470 4090 1500
rect 4380 1540 4470 1560
rect 4380 1500 4410 1540
rect 4450 1500 4470 1540
rect 4380 1460 4470 1500
rect 4380 1420 4410 1460
rect 4450 1420 4470 1460
rect 4380 1410 4470 1420
rect 3390 1310 4470 1410
use ring_vco  ring_vco_0
timestamp 1724224269
transform 1 0 900 0 1 3810
box -900 -3810 18620 2490
use sky130_fd_pr__res_generic_po_FARFDT  sky130_fd_pr__res_generic_po_FARFDT_0
timestamp 1724225640
transform 0 1 2865 -1 0 2550
box -40 -595 40 595
use sky130_fd_pr__res_generic_po_FARFDT  sky130_fd_pr__res_generic_po_FARFDT_1
timestamp 1724225640
transform 0 1 1525 -1 0 3170
box -40 -595 40 595
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 4488 0 -1 1762
box -38 -48 498 592
<< labels >>
rlabel metal1 3460 1570 3460 1570 1 VCCD
port 1 n
rlabel metal1 3460 1410 3460 1410 1 ENB
port 2 n
rlabel metal1 890 3210 890 3210 1 Anlg_in
port 4 n
<< end >>
