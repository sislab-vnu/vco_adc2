* NGSPICE file created from system.ext - technology: sky130A

.subckt count UP SetB DOWN Dout_buf GND VCCD
Xsky130_fd_sc_hd__dfstp_1_0 UP_buf Q2N SetBi GND GND VCCD VCCD Q1 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfstp_1_1 DWN_buf Q1_buf SetBi GND GND VCCD VCCD Q2 sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__inv_2_0 SetB GND GND VCCD VCCD SetBi sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_1 DOWN GND GND VCCD VCCD DWN_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_1 Q2 GND GND VCCD VCCD Q2N sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_2 Dout GND GND VCCD VCCD Dout_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_3 Q1 GND GND VCCD VCCD Q1_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_4 UP GND GND VCCD VCCD UP_buf sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__xor2_1_1 Q1 Q2 GND GND VCCD VCCD Dout sky130_fd_sc_hd__xor2_1
.ends

.subckt dco_freq clk clkDiv2 VNB VGND VPB VPWR
Xsky130_fd_sc_hd__buf_4_0 Q_N VGND VNB VPB VPWR Q_N_buf sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__inv_4_0 clk VGND VNB VPB VPWR clkinv sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__dfxtp_1_0 clkinv Q_N_buf VGND VNB VPB VPWR D sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxbp_2_0 clk D VGND VNB VPB VPWR clkDiv2 Q_N sky130_fd_sc_hd__dfxbp_2
.ends

.subckt dco_aux_inv VPWR VCCA A Y GND VGND
X0 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1
X1 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=1.2 ps=6.8 w=3 l=1
.ends

.subckt dco_main_inv VPWR VCCA Y GND VGND A
X0 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=1 M=2
X1 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=1 M=2
.ends

.subckt dco_cc_inv outp inp inn outn VCCA VGND VPWR GND
Xdco_aux_inv_0 VPWR VCCA outp outn GND VGND dco_aux_inv
Xdco_aux_inv_1 VPWR VCCA outn outp GND VGND dco_aux_inv
Xdco_main_inv_0 VPWR VCCA outp GND VGND inp dco_main_inv
Xdco_main_inv_1 VPWR VCCA outn GND VGND inn dco_main_inv
.ends

.subckt dco_ring_osc p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4] VGND p[0] VPWR
+ GND VCCA
Xdco_cc_inv_0 p[0] p[4] pn[4] pn[0] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_1 p[1] p[0] pn[0] pn[1] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_2 p[2] p[1] pn[1] pn[2] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_3 p[4] p[3] pn[3] pn[4] VCCA VGND VPWR GND dco_cc_inv
Xdco_cc_inv_4 p[3] p[2] pn[2] pn[3] VCCA VGND VPWR GND dco_cc_inv
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_RSCMUS a_n35_n1272# a_n35_840# a_n165_n1402#
X0 a_n35_840# a_n35_n1272# a_n165_n1402# sky130_fd_pr__res_xhigh_po_0p35 l=8.56
.ends

.subckt dco_idac Dctrl Vbs1 Vbs2 Vbs3 Vbs4 Isup VCCD VCCA GND
Xsky130_fd_sc_hd__buf_2_0 Dctrl GND GND VCCD VCCD G_M7 sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__inv_2_0 G_M7 GND GND VCCD VCCD G_M5 sky130_fd_sc_hd__inv_2
Xsky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0 GND D_M7 GND sky130_fd_pr__res_xhigh_po_0p35_RSCMUS
X0 Isup G_M7 D1_M4 GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X1 B_M2 Vbs1 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X2 D1_M4 Vbs4 D1_M3 D1_M3 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X3 D_M7 G_M5 D1_M4 GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5 M=2
X4 Isup G_M5 D1_M4 D1_M4 sky130_fd_pr__pfet_01v8_hvt ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.5 M=2
X5 D1_M3 Vbs3 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.2 as=0.72 ps=4.4 w=1.8 l=0.5 M=3
X6 Isup Vbs2 B_M2 B_M2 sky130_fd_pr__pfet_01v8_hvt ad=0.72 pd=4.4 as=0.72 ps=4.4 w=1.8 l=0.5
X7 D1_M4 G_M7 D_M7 D1_M4 sky130_fd_pr__pfet_01v8_hvt ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.5 M=2
.ends

.subckt dco VCCA Dctrl ENB Vbs_12 Vbs_34 pha_DCO GND Isup VCCD
Xdco_freq_0 pha_ro ro_div2 GND GND VCCD VCCD dco_freq
Xdco_freq_1 ro_div2 pha_DCO GND GND VCCD VCCD dco_freq
Xsky130_fd_sc_hd__buf_2_0 p_osc GND GND VCCD VCCD pha_ro sky130_fd_sc_hd__buf_2
Xdco_ring_osc_0 dco_ring_osc_0/p[1] dco_ring_osc_0/p[2] dco_ring_osc_0/p[3] p_osc
+ dco_ring_osc_0/pn[0] dco_ring_osc_0/pn[1] dco_ring_osc_0/pn[2] dco_ring_osc_0/pn[3]
+ dco_ring_osc_0/pn[4] GND dco_ring_osc_0/p[0] Isup GND Isup dco_ring_osc
Xdco_idac_0 Dctrl Vbs_12 Vbs_12 Vbs_34 Vbs_34 Isup VCCD VCCA GND dco_idac
Xsky130_fd_sc_hd__einvp_1_0 VCCD ENB GND GND VCCD VCCD dco_ring_osc_0/pn[4] sky130_fd_sc_hd__einvp_1
.ends

.subckt qz CLK Dout FBack D GND VCCD
Xsky130_fd_sc_hd__dlygate4sd3_1_0 CLK GND GND VCCD VCCD DL1 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_1 DL1 GND GND VCCD VCCD DL2 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__inv_2_0 FBack_inv GND GND VCCD VCCD FBack sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__buf_2_0 D GND GND VCCD VCCD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dlygate4sd3_1_2 DL2 GND GND VCCD VCCD DL3 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_3 DL3 GND GND VCCD VCCD DL4 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_4 DL4 GND GND VCCD VCCD DL5 sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__dlygate4sd3_1_5 DL5 GND GND VCCD VCCD CLK_dly sky130_fd_sc_hd__dlygate4sd3_1
Xsky130_fd_sc_hd__nand2_1_0 CLK_dly Dout GND GND VCCD VCCD FBack_inv sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfxtp_1_0 CLK sky130_fd_sc_hd__buf_2_0/X GND GND VCCD VCCD Dout
+ sky130_fd_sc_hd__dfxtp_1
.ends

.subckt sky130_fd_pr__res_generic_po_DKCPUZ a_n48_200# a_n48_n630#
R0 a_n48_200# a_n48_n630# sky130_fd_pr__res_generic_po w=0.48 l=2
.ends

.subckt mag_vco_main_inv A VPWR VGND Y VCCA GND
X0 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt mag_vco_aux_inv A VPWR VGND Y VCCA GND
X0 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt mag_vco_cc_inv inp inn VPWR VGND outp outn VCCA GND
Xmag_vco_main_inv_0 inp VPWR VGND outp VCCA GND mag_vco_main_inv
Xmag_vco_main_inv_1 inn VPWR VGND outn VCCA GND mag_vco_main_inv
Xmag_vco_aux_inv_0 outp VPWR VGND outn VCCA GND mag_vco_aux_inv
Xmag_vco_aux_inv_1 outn VPWR VGND outp VCCA GND mag_vco_aux_inv
.ends

.subckt mag_vco_ring_vco VGND p[0] p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4]
+ mag_vco_cc_inv_4/VCCA VSUBS VPWR
Xmag_vco_cc_inv_0 p[4] pn[4] VPWR VGND p[0] pn[0] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_1 p[0] pn[0] VPWR VGND p[1] pn[1] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_2 p[1] pn[1] VPWR VGND p[2] pn[2] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_3 p[3] pn[3] VPWR VGND p[4] pn[4] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_4 p[2] pn[2] VPWR VGND p[3] pn[3] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
.ends

.subckt vco VCCD ENB p[4] Anlg_in GND VCCA VPWR
Xsky130_fd_pr__res_generic_po_DKCPUZ_0 Anlg_in mag_vco_ring_vco_0/VGND sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_pr__res_generic_po_DKCPUZ_1 mag_vco_ring_vco_0/VGND GND sky130_fd_pr__res_generic_po_DKCPUZ
Xmag_vco_ring_vco_0 mag_vco_ring_vco_0/VGND mag_vco_ring_vco_0/p[0] mag_vco_ring_vco_0/p[1]
+ mag_vco_ring_vco_0/p[2] mag_vco_ring_vco_0/p[3] p[4] mag_vco_ring_vco_0/pn[0] mag_vco_ring_vco_0/pn[1]
+ mag_vco_ring_vco_0/pn[2] mag_vco_ring_vco_0/pn[3] mag_vco_ring_vco_0/pn[4] VCCA
+ GND VPWR mag_vco_ring_vco
Xsky130_fd_sc_hd__einvp_1_0 VCCD ENB GND GND VCCD VCCD mag_vco_ring_vco_0/pn[4] sky130_fd_sc_hd__einvp_1
.ends

.subckt system Dout CLK Anlg_in VCCD ENB GND Vbs_12 VCCA Vbs_34
Xcount_0 vco_0/p[4] ENB qz_0/FBack D1 GND VCCD count
Xdco_0 VCCA D1 ENB Vbs_12 Vbs_34 p_dco GND dco_0/Isup VCCD dco
Xcount_1 p_dco ENB qz_0/FBack qz_0/D GND VCCD count
Xqz_0 CLK Dout qz_0/FBack qz_0/D GND VCCD qz
Xvco_0 VCCD ENB vco_0/p[4] Anlg_in GND VCCA VCCA vco
.ends

