** sch_path: /home/toind/work/vco_adc2/xschem/lib_dco/dco_idac.sch
.subckt dco_idac VCCA Dctrl Vbs1 Vbs2 Vbs3 Vbs4 Isup
*.PININFO Vbs3:I Vbs4:I Vbs1:I Vbs2:I Isup:O Dctrl:I
x1 open GND GND VCCD VCCD lock sky130_fd_sc_hd__inv_2
XM1 note_12 Vbs1 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt L="L_br1" W="W_br1" nf=1 m=1
XM2 Isup Vbs2 note_12 note_12 sky130_fd_pr__pfet_01v8_hvt L="L_br1" W="W_br1" nf=1 m=1
x2 Dctrl GND GND VCCD VCCD open sky130_fd_sc_hd__buf_2
XM3 note_34 Vbs3 VCCA VCCA sky130_fd_pr__pfet_01v8_hvt L=L_br2 W="3*W_br2" nf=3 m=1
XM4 add_pwr Vbs4 note_34 note_34 sky130_fd_pr__pfet_01v8_hvt L=L_br2 W="3*W_br2" nf=3 m=1
XM5 Isup lock add_pwr add_pwr sky130_fd_pr__pfet_01v8_hvt L=Lp_lk W="2*Wp_lk" nf=2 m=1
XM6 add_pwr open Isup Isup sky130_fd_pr__nfet_01v8 L=Ln_lk W="2*Wn_lk" nf=2 m=1
XM7 input_R open add_pwr add_pwr sky130_fd_pr__pfet_01v8_hvt L=Lp_lk W="2*Wp_lk" nf=2 m=1
XM8 add_pwr lock input_R input_R sky130_fd_pr__nfet_01v8 L=Ln_lk W="2*Wn_lk" nf=2 m=1
XR2 GND input_R GND sky130_fd_pr__res_xhigh_po_0p35 L=8.562 mult=1 m=1
.ends
.GLOBAL GND
.end
