magic
tech sky130A
timestamp 1729593089
<< locali >>
rect 2980 1375 3090 1415
rect 5980 1375 6090 1415
rect 8880 1375 10020 1415
rect 2980 150 3090 190
rect 3095 -690 3145 170
rect 5980 150 6090 190
rect 5910 -725 6020 -685
rect 8860 -695 8910 180
rect 9920 -1910 10020 1375
rect 5910 -1950 6020 -1910
rect 8825 -1950 10020 -1910
<< metal1 >>
rect 20 1515 120 1565
rect 1955 1515 3055 1565
rect 4935 1515 6110 1565
rect 8005 1515 9765 1565
rect -300 1075 0 1125
rect 2980 1075 3090 1125
rect 5980 1075 6090 1125
rect 9000 1075 9490 1125
rect -300 -1610 -250 1075
rect -150 440 0 490
rect 2980 440 3090 490
rect 5980 440 6090 490
rect 9000 440 9200 490
rect -150 -975 -100 440
rect 2025 0 3050 50
rect 3900 -540 3950 25
rect 5035 0 6045 50
rect 5930 -585 6955 -535
rect 8050 -570 8100 50
rect 9100 -975 9200 440
rect -150 -1025 3000 -975
rect 5910 -1025 6020 -975
rect 9000 -1025 9200 -975
rect 9390 -1610 9490 1075
rect -300 -1660 3000 -1610
rect 5910 -1660 6020 -1610
rect 9000 -1660 9490 -1610
rect 9665 -2050 9765 1515
rect 5875 -2100 6925 -2050
rect 8875 -2100 9765 -2050
use vco_cc_inv  vco_cc_inv_0
timestamp 1729593089
transform 1 0 130 0 1 150
box -130 -150 2870 1415
use vco_cc_inv  vco_cc_inv_1
timestamp 1729593089
transform 1 0 3130 0 1 150
box -130 -150 2870 1415
use vco_cc_inv  vco_cc_inv_2
timestamp 1729593089
transform 1 0 6130 0 1 150
box -130 -150 2870 1415
use vco_cc_inv  vco_cc_inv_3
timestamp 1729593089
transform -1 0 5870 0 -1 -685
box -130 -150 2870 1415
use vco_cc_inv  vco_cc_inv_4
timestamp 1729593089
transform -1 0 8870 0 -1 -685
box -130 -150 2870 1415
<< labels >>
rlabel locali s 3095 -255 3095 -255 4 VGND
rlabel locali s 2990 1415 2990 1415 4 VPWR
rlabel metal1 s 3040 1125 3040 1125 4 p[0]
rlabel metal1 s 6035 1125 6035 1125 4 p[1]
rlabel metal1 s 9125 1125 9125 1125 4 p[2]
rlabel metal1 s 5965 -1610 5965 -1610 4 p[3]
rlabel metal1 s 2945 -1610 2945 -1610 4 p[4]
rlabel metal1 s 3035 490 3035 490 4 pn[0]
rlabel metal1 s 6035 490 6035 490 4 pn[1]
rlabel metal1 s 9095 490 9095 490 4 pn[2]
rlabel metal1 s 5960 -975 5960 -975 4 pn[3]
rlabel metal1 s 2940 -975 2940 -975 4 pn[4]
rlabel metal1 s 30 1565 30 1565 4 VCCA
rlabel metal1 s 3950 -500 3950 -500 4 GND
<< end >>
