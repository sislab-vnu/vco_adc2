* NGSPICE file created from mag_vco_ring_vco.ext - technology: sky130A

.subckt mag_vco_main_inv A VPWR VGND Y VCCA GND
X0 VPWR A Y VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt mag_vco_aux_inv A VPWR VGND Y VCCA GND
X0 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt mag_vco_cc_inv inp inn VPWR VGND outp outn VCCA GND
Xmag_vco_main_inv_0 inp VPWR VGND outp VCCA GND mag_vco_main_inv
Xmag_vco_main_inv_1 inn VPWR VGND outn VCCA GND mag_vco_main_inv
Xmag_vco_aux_inv_0 outp VPWR VGND outn VCCA GND mag_vco_aux_inv
Xmag_vco_aux_inv_1 outn VPWR VGND outp VCCA GND mag_vco_aux_inv
.ends

.subckt mag_vco_ring_vco VGND VPWR p[0] p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3]
+ pn[4]
Xmag_vco_cc_inv_0 p[4] pn[4] VPWR VGND p[0] pn[0] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_2 p[1] pn[1] VPWR VGND p[2] pn[2] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_1 p[0] pn[0] VPWR VGND p[1] pn[1] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_3 p[3] pn[3] VPWR VGND p[4] pn[4] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
Xmag_vco_cc_inv_4 p[2] pn[2] VPWR VGND p[3] pn[3] mag_vco_cc_inv_4/VCCA VSUBS mag_vco_cc_inv
.ends

