magic
tech sky130A
magscale 1 2
timestamp 1727091651
<< locali >>
rect -3015 4470 2150 4580
rect -3060 4110 3220 4150
rect -3060 4070 3130 4110
rect 3170 4070 3220 4110
rect -3060 4050 3220 4070
rect -4470 3590 2990 3650
rect -4470 -1750 -4410 3590
rect -4470 -1830 1430 -1750
rect -4470 -3890 -4410 -1830
rect -3300 -2860 -3200 -2830
rect -3300 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3300 -2920 -3200 -2900
rect 1350 -3350 1430 -1830
rect 15700 -1800 15770 -1260
rect 15700 -1840 15720 -1800
rect 15760 -1840 15770 -1800
rect 15700 -1860 15770 -1840
rect 19560 -2490 21710 -2480
rect 19560 -2530 19580 -2490
rect 19620 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 19560 -2550 21710 -2530
rect 18400 -3070 18470 -2660
rect 1350 -3370 5570 -3350
rect 1350 -3410 5520 -3370
rect 5560 -3410 5570 -3370
rect 1350 -3430 5570 -3410
rect -4470 -3930 -4460 -3890
rect -4420 -3930 -4410 -3890
rect -4470 -11680 -4410 -3930
rect 390 -4850 570 -4820
rect 390 -4890 500 -4850
rect 540 -4890 570 -4850
rect 390 -4920 570 -4890
rect 14840 -7240 15030 -7200
rect 14840 -7270 15490 -7240
rect 14840 -7320 14910 -7270
rect 14960 -7320 15490 -7270
rect 14840 -7380 15030 -7320
rect 15280 -8300 15380 -8270
rect 15280 -8340 15310 -8300
rect 15350 -8340 15380 -8300
rect 15280 -11680 15380 -8340
rect 19080 -9260 19180 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 19180 -9260
rect 19080 -9330 19180 -9300
rect -4470 -11780 15380 -11680
<< viali >>
rect 540 7650 580 7690
rect 1630 7650 1670 7690
rect 2720 7650 2760 7690
rect 4640 7650 4680 7690
rect 6540 7650 6580 7690
rect 7630 7650 7670 7690
rect 8720 7650 8760 7690
rect 10640 7650 10680 7690
rect 12540 7650 12580 7690
rect 13630 7650 13670 7690
rect 14720 7650 14760 7690
rect 17420 7650 17460 7690
rect 3130 4070 3170 4110
rect 6400 1000 6440 1040
rect 7490 1000 7530 1040
rect 8580 1000 8620 1040
rect 10480 1000 10520 1040
rect 12400 1000 12440 1040
rect 13490 1000 13530 1040
rect 14580 1000 14620 1040
rect 16480 1000 16520 1040
rect 17420 1000 17460 1040
rect 740 -2610 780 -2570
rect -3270 -2900 -3230 -2860
rect 15720 -1840 15760 -1800
rect 19580 -2530 19620 -2490
rect 21650 -2530 21690 -2490
rect 5520 -3410 5560 -3370
rect -4460 -3930 -4420 -3890
rect 500 -4890 540 -4850
rect 14910 -7320 14960 -7270
rect 15310 -8340 15350 -8300
rect 19110 -9300 19150 -9260
<< metal1 >>
rect -2080 7910 -1310 8010
rect -3390 1560 -1760 1660
rect -3390 -2830 -3300 1560
rect 14930 -1600 15640 -1500
rect 730 -2560 1240 -2550
rect 730 -2570 780 -2560
rect 730 -2610 740 -2570
rect 730 -2620 780 -2610
rect 840 -2620 1240 -2560
rect 730 -2630 1240 -2620
rect -3390 -2860 -3200 -2830
rect -3390 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3390 -2920 -3200 -2900
rect 5500 -3370 5570 -3350
rect 5500 -3410 5520 -3370
rect 5560 -3410 5570 -3370
rect 5500 -3430 5570 -3410
rect -4470 -3890 -3160 -3870
rect -4470 -3930 -4460 -3890
rect -4420 -3930 -3160 -3890
rect -4470 -3950 -3160 -3930
rect -70 -3970 60 -3960
rect -70 -4030 -10 -3970
rect 50 -4030 60 -3970
rect -70 -4040 60 -4030
rect 470 -4850 570 -4820
rect 470 -4890 500 -4850
rect 540 -4890 570 -4850
rect 470 -12490 570 -4890
rect 14930 -5475 15030 -1600
rect 19560 -2490 19640 -2470
rect 19560 -2530 19580 -2490
rect 19620 -2530 19640 -2490
rect 19560 -2550 19640 -2530
rect 21610 -2490 21710 -2480
rect 21610 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 15480 -2640 15800 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2690 15800 -2640
rect 15560 -2700 15580 -2690
rect 15480 -2720 15580 -2700
rect 10995 -5565 15720 -5475
rect 15630 -6940 15720 -5565
rect 14840 -7260 15030 -7200
rect 14840 -7330 14900 -7260
rect 14970 -7330 15030 -7260
rect 14840 -7380 15030 -7330
rect 15280 -8286 15380 -8270
rect 15280 -8300 15570 -8286
rect 15280 -8340 15310 -8300
rect 15350 -8340 15570 -8300
rect 15280 -8356 15570 -8340
rect 15280 -8370 15380 -8356
rect 18700 -8376 18800 -8360
rect 18540 -8380 18800 -8376
rect 18540 -8440 18720 -8380
rect 18780 -8440 18800 -8380
rect 18540 -8446 18800 -8440
rect 18700 -8460 18800 -8446
rect 21610 -9230 21710 -2530
rect 19080 -9260 21710 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 21710 -9260
rect 19080 -9330 21710 -9300
rect 21610 -12490 21710 -9330
rect 470 -12590 21710 -12490
<< via1 >>
rect 780 -2620 840 -2560
rect -10 -4030 50 -3970
rect 15500 -2700 15560 -2640
rect 14900 -7270 14970 -7260
rect 14900 -7320 14910 -7270
rect 14910 -7320 14960 -7270
rect 14960 -7320 14970 -7270
rect 14900 -7330 14970 -7320
rect 3870 -8260 3930 -8200
rect 18720 -8440 18780 -8380
<< metal2 >>
rect 730 -2560 2000 -2550
rect 730 -2620 780 -2560
rect 840 -2620 2000 -2560
rect 730 -2630 2000 -2620
rect 15480 -2640 15580 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2700 15580 -2640
rect -20 -3970 1000 -3960
rect -20 -4030 -10 -3970
rect 50 -4030 1000 -3970
rect -20 -4040 1000 -4030
rect 920 -7670 1000 -4040
rect 15480 -6300 15580 -2700
rect 15480 -6400 19700 -6300
rect 14840 -7260 15030 -7200
rect 14840 -7330 14900 -7260
rect 14970 -7330 15030 -7260
rect 14840 -7380 15030 -7330
rect 920 -7750 3940 -7670
rect 3860 -8180 3940 -7750
rect 3850 -8200 3950 -8180
rect 3850 -8260 3870 -8200
rect 3930 -8260 3950 -8200
rect 3850 -8270 3950 -8260
rect 14869 -9240 14972 -7380
rect 19600 -8360 19700 -6400
rect 18700 -8380 19700 -8360
rect 18700 -8440 18720 -8380
rect 18780 -8440 19700 -8380
rect 18700 -8460 19700 -8440
rect 14330 -9340 14972 -9240
rect 14869 -9341 14972 -9340
use count  count_0 ../count
timestamp 1727087206
transform 1 0 -2340 0 1 -2076
box -880 -3154 3140 -440
use count  count_1
timestamp 1727087206
transform 1 0 16330 0 1 -6486
box -880 -3154 3140 -440
use dco  dco_0 ../dco
timestamp 1727083693
transform 1 0 2620 0 1 -6850
box -720 -4280 11940 6160
use qz  qz_0 ../quantizer
timestamp 1727065578
transform 1 0 15260 0 1 -2230
box 190 -710 5890 730
use vco  vco_0 ../vco_v3
timestamp 1725958133
transform 1 0 -2020 0 1 680
box 0 0 19930 7330
<< labels >>
flabel space -2990 4650 -2990 4650 0 FreeSans 1600 0 0 0 1
flabel space -3040 4200 -3040 4200 0 FreeSans 1600 0 0 0 2
flabel space -3050 3680 -3050 3680 0 FreeSans 1600 0 0 0 3
flabel space -2020 8090 -2020 8090 0 FreeSans 1600 0 0 0 4
flabel space -3330 1750 -3330 1750 0 FreeSans 1600 0 0 0 5
flabel space -3980 -3760 -3970 -3760 0 FreeSans 1600 0 0 0 6
flabel space 1010 -3860 1010 -3860 0 FreeSans 1600 0 0 0 7
flabel space 5290 -3500 5290 -3500 0 FreeSans 1600 0 0 0 8
flabel space 5200 -5820 5200 -5820 0 FreeSans 1600 0 0 0 9
flabel space 6660 -6200 6660 -6200 0 FreeSans 1600 0 0 0 10
flabel space 4400 -660 4400 -660 0 FreeSans 1600 0 0 0 11
flabel space 1910 -510 1910 -510 0 FreeSans 1600 0 0 0 12
flabel space 15010 -7110 15010 -7110 0 FreeSans 1600 0 0 0 13
flabel space 15190 -8110 15190 -8110 0 FreeSans 1600 0 0 0 14
flabel space 18880 -8310 18880 -8310 0 FreeSans 1600 0 0 0 15
flabel space 15710 -1220 15710 -1220 0 FreeSans 1600 0 0 0 16
flabel space 18370 -3200 18370 -3200 0 FreeSans 1600 0 0 0 17
<< end >>
