magic
tech sky130A
timestamp 1723792769
<< nwell >>
rect 4065 105 4130 265
rect -222 -405 -136 -403
rect -222 -566 -117 -405
rect 1101 -580 1264 -359
rect 1100 -710 1360 -580
rect 2234 -710 2560 -580
rect 2234 -1150 2314 -710
rect 1456 -1476 1551 -1315
rect 1770 -1475 1990 -1315
<< pwell >>
rect 4045 -15 4130 75
rect -167 -686 -100 -618
rect 1444 -1060 1545 -820
rect 1780 -1060 1880 -820
rect 1480 -1596 1570 -1527
rect 1750 -1596 2012 -1505
<< psubdiff >>
rect 4075 40 4105 55
rect 4075 20 4080 40
rect 4100 20 4105 40
rect 4075 5 4105 20
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
rect 1471 -954 1501 -937
rect 1471 -971 1478 -954
rect 1495 -971 1501 -954
rect 1471 -987 1501 -971
rect 1499 -1553 1529 -1536
rect 1499 -1570 1506 -1553
rect 1523 -1570 1529 -1553
rect 1499 -1586 1529 -1570
<< nsubdiff >>
rect 4075 165 4105 180
rect 4075 145 4080 165
rect 4100 145 4105 165
rect 4075 130 4105 145
rect -165 -484 -135 -467
rect -165 -501 -158 -484
rect -141 -501 -135 -484
rect -165 -517 -135 -501
rect 1147 -517 1177 -501
rect 1147 -534 1154 -517
rect 1171 -534 1177 -517
rect 1147 -551 1177 -534
rect 2401 -638 2431 -620
rect 2401 -655 2408 -638
rect 2425 -655 2431 -638
rect 2401 -670 2431 -655
rect 1492 -1382 1522 -1365
rect 1492 -1399 1498 -1382
rect 1515 -1399 1522 -1382
rect 1492 -1415 1522 -1399
<< psubdiffcont >>
rect 4080 20 4100 40
rect -148 -661 -130 -644
rect 1478 -971 1495 -954
rect 1506 -1570 1523 -1553
<< nsubdiffcont >>
rect 4080 145 4100 165
rect -158 -501 -141 -484
rect 1154 -534 1171 -517
rect 2408 -655 2425 -638
rect 1498 -1399 1515 -1382
<< locali >>
rect 4075 165 4105 180
rect 4075 145 4080 165
rect 4100 145 4105 165
rect 4075 130 4105 145
rect 3995 84 4207 105
rect 200 -450 270 50
rect 4075 40 4105 55
rect 4075 20 4080 40
rect 4100 20 4105 40
rect 4075 5 4105 20
rect 4167 -222 4207 84
rect 4167 -239 4179 -222
rect 4196 -239 4207 -222
rect 4167 -246 4207 -239
rect -165 -484 -135 -467
rect 120 -480 270 -450
rect -165 -501 -158 -484
rect -141 -501 -135 -484
rect -165 -517 -135 -501
rect 1147 -517 1177 -501
rect 1147 -534 1154 -517
rect 1171 -534 1177 -517
rect 1147 -551 1177 -534
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
rect 2401 -638 2431 -620
rect 2401 -655 2408 -638
rect 2425 -655 2431 -638
rect 2401 -670 2431 -655
rect 1471 -954 1501 -937
rect 1471 -971 1478 -954
rect 1495 -971 1501 -954
rect 1471 -987 1501 -971
rect 1492 -1382 1522 -1365
rect 1492 -1399 1498 -1382
rect 1515 -1399 1522 -1382
rect 1492 -1415 1522 -1399
rect 1499 -1553 1529 -1536
rect 1499 -1570 1506 -1553
rect 1523 -1570 1529 -1553
rect 1499 -1586 1529 -1570
<< viali >>
rect 4080 145 4100 165
rect 3883 82 3900 99
rect 4080 20 4100 40
rect 4179 -239 4196 -222
rect 1154 -534 1171 -517
rect -70 -590 -50 -570
rect 99 -589 116 -572
rect -148 -661 -130 -644
rect 2408 -655 2425 -638
rect 4135 -719 4152 -702
rect 1478 -971 1495 -954
rect 1498 -1399 1515 -1382
rect 4135 -1525 4152 -1508
rect 1506 -1570 1523 -1553
<< metal1 >>
rect 4075 165 4105 180
rect 3416 109 3450 150
rect 4075 145 4080 165
rect 4100 145 4105 165
rect 4075 130 4105 145
rect 3416 99 3908 109
rect 3416 82 3883 99
rect 3900 82 3908 99
rect 3416 73 3908 82
rect 4075 40 4105 55
rect 4075 20 4080 40
rect 4100 20 4105 40
rect 4075 5 4105 20
rect 1370 -200 1630 -160
rect 2040 -200 2290 -160
rect -165 -517 -135 -467
rect 1147 -517 1177 -501
rect 1147 -534 1154 -517
rect 1171 -534 1177 -517
rect 1147 -551 1177 -534
rect -90 -570 -47 -555
rect -140 -590 -70 -570
rect -50 -590 -47 -570
rect -140 -600 -47 -590
rect 96 -571 121 -558
rect 96 -572 169 -571
rect 96 -589 99 -572
rect 116 -589 169 -572
rect 96 -605 121 -589
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
rect 2401 -638 2431 -620
rect 2401 -655 2408 -638
rect 2425 -655 2431 -638
rect 2401 -670 2431 -655
rect 1471 -954 1501 -937
rect 1471 -971 1478 -954
rect 1495 -971 1501 -954
rect 1471 -987 1501 -971
rect 2685 -1230 2735 -80
rect 4127 -702 4160 -693
rect 4127 -719 4135 -702
rect 4152 -719 4160 -702
rect 4127 -754 4160 -719
rect 3813 -783 4160 -754
rect 3813 -1016 3842 -783
rect 2643 -1270 2735 -1230
rect 1492 -1382 1522 -1365
rect 1492 -1399 1498 -1382
rect 1515 -1399 1522 -1382
rect 1492 -1415 1522 -1399
rect 1223 -1508 1482 -1471
rect 4127 -1508 4160 -1497
rect 4127 -1525 4135 -1508
rect 4152 -1525 4160 -1508
rect 1499 -1553 1529 -1536
rect 1499 -1570 1506 -1553
rect 1523 -1570 1529 -1553
rect 4127 -1554 4160 -1525
rect 1499 -1586 1529 -1570
rect 3815 -1584 4160 -1554
rect 3815 -1773 3845 -1584
use div_d  div_d_0
timestamp 1723787705
transform 1 0 4271 0 1 -1262
box -921 312 740 1046
use div_d  div_d_1
timestamp 1723787705
transform 1 0 4271 0 1 -2062
box -921 312 740 1046
use idac_p  idac_p_0
timestamp 1723776395
transform 1 0 1480 0 1 -580
box -380 -1170 1163 420
use ring_osc_d  ring_osc_d_0
timestamp 1723780164
transform 1 0 180 0 1 810
box -280 -900 5060 750
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3864 0 1 -26
box -19 -24 203 296
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -101 0 1 -696
box -19 -24 249 296
<< end >>
