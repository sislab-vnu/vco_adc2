VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc2
  CLASS BLOCK ;
  FOREIGN vco_adc2 ;
  ORIGIN 37.950 320.620 ;
  SIZE 171.570 BY 505.310 ;
  PIN vbias_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 38.900 -25.650 39.200 -25.150 ;
        RECT 53.450 -25.700 53.950 -25.200 ;
      LAYER met1 ;
        RECT 32.700 -22.500 33.700 -22.300 ;
        RECT 32.700 -23.000 53.950 -22.500 ;
        RECT 32.700 -23.300 33.700 -23.000 ;
        RECT 40.250 -25.150 40.750 -23.000 ;
        RECT 38.700 -25.650 40.750 -25.150 ;
        RECT 53.450 -25.700 53.950 -23.000 ;
      LAYER met2 ;
        RECT 22.650 -23.300 33.700 -22.300 ;
        RECT 22.650 -318.100 24.650 -23.300 ;
        RECT 22.650 -320.100 133.350 -318.100 ;
      LAYER met3 ;
        RECT 125.460 -320.620 133.620 -317.900 ;
    END
  END vbias_12
  PIN vbias_34
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER li1 ;
        RECT 42.650 -25.650 43.650 -25.150 ;
        RECT 47.950 -25.650 50.250 -25.150 ;
      LAYER met1 ;
        RECT 45.500 -25.150 46.500 -24.650 ;
        RECT 42.450 -25.650 50.250 -25.150 ;
      LAYER met2 ;
        RECT 45.500 -24.450 58.400 -23.450 ;
        RECT 45.500 -25.650 46.500 -24.450 ;
        RECT 57.400 -52.800 58.400 -24.450 ;
        RECT 57.400 -54.850 132.150 -52.800 ;
      LAYER met3 ;
        RECT 124.440 -55.420 132.600 -52.020 ;
    END
  END vbias_34
  PIN analog_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.000 24.600 34.500 24.700 ;
        RECT 29.185 24.280 34.500 24.600 ;
        RECT 31.000 24.000 34.500 24.280 ;
      LAYER met1 ;
        RECT 34.500 24.700 35.700 25.000 ;
        RECT 29.125 24.250 31.230 24.630 ;
        RECT 33.500 24.000 35.700 24.700 ;
      LAYER met2 ;
        RECT 86.710 176.600 88.550 184.690 ;
        RECT 86.710 174.600 124.950 176.600 ;
        RECT 86.710 174.570 88.550 174.600 ;
        RECT 122.950 25.000 124.950 174.600 ;
        RECT 34.500 24.000 124.950 25.000 ;
    END
  END analog_in
  PIN enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.437000 ;
    PORT
      LAYER li1 ;
        RECT -14.150 20.050 15.300 20.250 ;
        RECT 15.625 20.050 16.085 20.115 ;
        RECT -14.150 19.750 16.085 20.050 ;
        RECT -14.150 19.250 -13.650 19.750 ;
        RECT 11.600 4.650 12.100 19.750 ;
        RECT 15.625 19.385 16.085 19.750 ;
        RECT 11.600 4.150 30.150 4.650 ;
        RECT 29.650 -5.900 30.150 4.150 ;
        RECT 29.650 -6.400 35.200 -5.900 ;
        RECT -8.955 -7.575 -8.625 -7.325 ;
        RECT 34.700 -8.450 35.200 -6.400 ;
        RECT 34.700 -8.950 41.450 -8.450 ;
        RECT 42.525 -8.765 42.985 -8.035 ;
        RECT -14.150 -38.850 -13.650 -38.350 ;
        RECT -14.150 -39.350 -9.450 -38.850 ;
        RECT -8.955 -39.225 -8.625 -38.975 ;
      LAYER met1 ;
        RECT -14.150 -7.150 -13.150 20.250 ;
        RECT 13.550 19.750 15.300 20.250 ;
        RECT -14.150 -7.280 -10.000 -7.150 ;
        RECT -14.150 -7.630 -8.600 -7.280 ;
        RECT -14.150 -7.650 -10.000 -7.630 ;
        RECT -14.150 -39.350 -13.150 -7.650 ;
        RECT 39.950 -8.500 41.450 -8.450 ;
        RECT 42.500 -8.500 43.000 -8.250 ;
        RECT 39.950 -8.800 43.000 -8.500 ;
        RECT 39.950 -8.950 41.450 -8.800 ;
        RECT -10.500 -38.930 -9.450 -38.850 ;
        RECT -10.500 -39.280 -8.600 -38.930 ;
        RECT -10.500 -39.350 -9.450 -39.280 ;
      LAYER met2 ;
        RECT -37.600 17.250 -13.150 19.250 ;
        RECT -37.600 -88.850 -35.600 17.250 ;
        RECT -14.150 16.250 -13.150 17.250 ;
        RECT -37.950 -94.830 -35.190 -88.850 ;
    END
  END enable_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER li1 ;
        RECT -7.325 -21.405 -6.635 -20.845 ;
        RECT -3.520 -25.485 -3.170 -24.835 ;
      LAYER met1 ;
        RECT -7.320 -20.950 -6.620 -20.830 ;
        RECT -8.850 -21.300 -6.620 -20.950 ;
        RECT -8.850 -22.950 -7.850 -21.300 ;
        RECT -7.320 -21.400 -6.620 -21.300 ;
        RECT -8.850 -23.300 -4.000 -22.950 ;
        RECT -4.350 -24.800 -4.000 -23.300 ;
        RECT -4.350 -24.840 -3.200 -24.800 ;
        RECT -4.350 -25.150 -3.190 -24.840 ;
        RECT -3.540 -25.490 -3.190 -25.150 ;
      LAYER met2 ;
        RECT -25.850 -18.800 -7.850 -17.800 ;
        RECT -25.850 -86.500 -23.850 -18.800 ;
        RECT -8.850 -23.300 -7.850 -18.800 ;
        RECT -25.850 -87.300 -16.900 -86.500 ;
        RECT -25.850 -88.500 -16.930 -87.300 ;
        RECT -19.690 -94.830 -16.930 -88.500 ;
    END
  END clk
  PIN quantizer_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 3.275 -24.885 3.605 -24.040 ;
        RECT 3.275 -24.965 3.665 -24.885 ;
        RECT 3.450 -25.015 3.665 -24.965 ;
        RECT 3.495 -25.150 3.665 -25.015 ;
        RECT 5.735 -25.150 6.070 -25.135 ;
        RECT 3.495 -25.400 6.070 -25.150 ;
        RECT 3.495 -25.595 3.665 -25.400 ;
        RECT 3.440 -25.635 3.665 -25.595 ;
        RECT 3.285 -25.720 3.665 -25.635 ;
        RECT 3.285 -26.155 3.615 -25.720 ;
        RECT 4.300 -29.350 5.300 -25.400 ;
        RECT 5.735 -25.405 6.070 -25.400 ;
      LAYER met1 ;
        RECT 4.300 -29.350 6.400 -28.350 ;
      LAYER met2 ;
        RECT 5.300 -29.350 16.150 -28.350 ;
        RECT 14.150 -88.850 16.150 -29.350 ;
        RECT 14.030 -94.830 16.790 -88.850 ;
    END
  END quantizer_out
  PIN VDDA
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -7.100 33.650 82.900 39.450 ;
        RECT 15.350 19.700 18.750 21.300 ;
        RECT 15.350 19.695 18.030 19.700 ;
        RECT 22.900 7.600 82.900 13.400 ;
        RECT -10.000 -2.180 7.750 -0.480 ;
        RECT -9.950 -5.740 -9.050 -5.680 ;
        RECT -9.950 -7.345 -7.490 -5.740 ;
        RECT 2.350 -6.210 3.350 -6.180 ;
        RECT -9.950 -7.380 -9.100 -7.345 ;
        RECT -1.240 -7.815 5.560 -6.210 ;
        RECT 2.350 -7.830 3.350 -7.815 ;
        RECT 41.400 -8.450 44.930 -6.850 ;
        RECT 42.250 -8.455 44.930 -8.450 ;
        RECT -6.650 -12.395 -5.800 -12.380 ;
        RECT 4.100 -12.395 5.900 -12.380 ;
        RECT -8.390 -14.000 7.890 -12.395 ;
        RECT -6.650 -14.030 -5.800 -14.000 ;
        RECT 4.100 -14.030 6.050 -14.000 ;
        RECT -7.400 -19.550 17.300 -19.500 ;
        RECT -7.600 -21.200 17.300 -19.550 ;
        RECT 59.850 -21.850 62.700 -20.250 ;
        RECT 59.850 -21.855 62.070 -21.850 ;
        RECT -6.450 -23.550 9.900 -23.500 ;
        RECT -7.600 -25.200 9.900 -23.550 ;
        RECT 65.550 -24.150 67.700 -24.100 ;
        RECT 37.400 -28.250 39.800 -25.650 ;
        RECT 41.150 -28.250 45.350 -25.650 ;
        RECT 65.550 -25.750 79.940 -24.150 ;
        RECT 67.600 -25.755 79.940 -25.750 ;
        RECT 70.200 -25.800 72.300 -25.755 ;
        RECT 64.550 -29.950 82.300 -28.350 ;
        RECT 65.400 -29.955 82.300 -29.950 ;
        RECT 68.500 -30.000 70.850 -29.955 ;
        RECT 80.800 -30.000 82.300 -29.955 ;
        RECT -10.000 -33.830 7.750 -32.130 ;
        RECT 32.545 -37.250 34.150 -35.100 ;
        RECT -9.950 -37.390 -9.050 -37.330 ;
        RECT -9.950 -38.995 -7.490 -37.390 ;
        RECT 2.350 -37.860 3.350 -37.830 ;
        RECT -9.950 -39.030 -9.100 -38.995 ;
        RECT -1.240 -39.465 5.560 -37.860 ;
        RECT 32.500 -38.400 34.150 -37.250 ;
        RECT 65.550 -35.850 67.700 -35.800 ;
        RECT 65.550 -37.450 79.940 -35.850 ;
        RECT 67.600 -37.455 79.940 -37.450 ;
        RECT 70.200 -37.500 72.300 -37.455 ;
        RECT 2.350 -39.480 3.350 -39.465 ;
        RECT 32.545 -40.160 34.150 -38.400 ;
        RECT 64.550 -41.650 82.300 -40.050 ;
        RECT 65.400 -41.655 82.300 -41.650 ;
        RECT 68.500 -41.700 70.850 -41.655 ;
        RECT 80.800 -41.700 82.300 -41.655 ;
        RECT -6.650 -44.045 -5.800 -44.030 ;
        RECT 4.100 -44.045 5.900 -44.030 ;
        RECT -8.390 -45.650 7.890 -44.045 ;
        RECT -6.650 -45.680 -5.800 -45.650 ;
        RECT 4.100 -45.680 6.050 -45.650 ;
      LAYER li1 ;
        RECT -6.900 39.950 93.100 40.350 ;
        RECT -6.900 38.600 -6.500 39.950 ;
        RECT -6.200 34.050 -5.800 39.950 ;
        RECT 1.900 34.050 2.300 39.950 ;
        RECT 2.600 39.050 3.000 39.950 ;
        RECT 3.300 39.050 3.700 39.950 ;
        RECT 2.600 38.600 3.700 39.050 ;
        RECT 8.050 39.050 8.450 39.950 ;
        RECT 8.750 39.050 9.150 39.950 ;
        RECT 8.050 38.600 9.150 39.050 ;
        RECT 13.500 38.600 13.900 39.950 ;
        RECT 3.300 34.050 3.700 38.600 ;
        RECT 8.750 34.050 9.150 38.600 ;
        RECT 14.200 34.050 14.600 39.950 ;
        RECT 22.300 34.050 22.700 39.950 ;
        RECT 23.100 38.600 23.500 39.950 ;
        RECT 23.800 34.050 24.200 39.950 ;
        RECT 31.900 34.050 32.300 39.950 ;
        RECT 32.600 39.050 33.000 39.950 ;
        RECT 33.300 39.050 33.700 39.950 ;
        RECT 32.600 38.600 33.700 39.050 ;
        RECT 38.050 39.050 38.450 39.950 ;
        RECT 38.750 39.050 39.150 39.950 ;
        RECT 38.050 38.600 39.150 39.050 ;
        RECT 43.500 38.600 43.900 39.950 ;
        RECT 33.300 34.050 33.700 38.600 ;
        RECT 38.750 34.050 39.150 38.600 ;
        RECT 44.200 34.050 44.600 39.950 ;
        RECT 52.300 34.050 52.700 39.950 ;
        RECT 53.100 38.600 53.500 39.950 ;
        RECT 53.800 34.050 54.200 39.950 ;
        RECT 61.900 34.050 62.300 39.950 ;
        RECT 62.600 39.050 63.000 39.950 ;
        RECT 63.300 39.050 63.700 39.950 ;
        RECT 62.600 38.600 63.700 39.050 ;
        RECT 68.050 39.050 68.450 39.950 ;
        RECT 68.750 39.050 69.150 39.950 ;
        RECT 68.050 38.600 69.150 39.050 ;
        RECT 73.500 38.600 73.900 39.950 ;
        RECT 63.300 34.050 63.700 38.600 ;
        RECT 68.750 34.050 69.150 38.600 ;
        RECT 74.200 34.050 74.600 39.950 ;
        RECT 82.300 34.050 82.700 39.950 ;
        RECT 15.540 21.025 17.840 21.195 ;
        RECT 16.055 20.625 16.990 21.025 ;
        RECT 17.515 20.050 17.755 20.345 ;
        RECT 18.100 20.250 18.500 20.750 ;
        RECT 17.515 19.550 17.950 20.050 ;
        RECT 17.515 19.365 17.755 19.550 ;
        RECT 19.150 7.100 19.650 20.050 ;
        RECT 23.100 7.100 23.500 13.000 ;
        RECT 31.200 7.100 31.600 13.000 ;
        RECT 36.650 8.450 37.050 13.000 ;
        RECT 42.100 8.450 42.500 13.000 ;
        RECT 31.900 7.100 32.300 8.450 ;
        RECT 36.650 8.000 37.750 8.450 ;
        RECT 36.650 7.100 37.050 8.000 ;
        RECT 37.350 7.100 37.750 8.000 ;
        RECT 42.100 8.000 43.200 8.450 ;
        RECT 42.100 7.100 42.500 8.000 ;
        RECT 42.800 7.100 43.200 8.000 ;
        RECT 43.500 7.100 43.900 13.000 ;
        RECT 51.600 7.100 52.000 13.000 ;
        RECT 52.300 7.100 52.700 8.450 ;
        RECT 53.100 7.100 53.500 13.000 ;
        RECT 61.200 7.100 61.600 13.000 ;
        RECT 66.650 8.450 67.050 13.000 ;
        RECT 72.100 8.450 72.500 13.000 ;
        RECT 61.900 7.100 62.300 8.450 ;
        RECT 66.650 8.000 67.750 8.450 ;
        RECT 66.650 7.100 67.050 8.000 ;
        RECT 67.350 7.100 67.750 8.000 ;
        RECT 72.100 8.000 73.200 8.450 ;
        RECT 72.100 7.100 72.500 8.000 ;
        RECT 72.800 7.100 73.200 8.000 ;
        RECT 73.500 7.100 73.900 13.000 ;
        RECT 81.600 7.100 82.000 13.000 ;
        RECT 82.300 7.100 82.700 8.450 ;
        RECT 92.100 7.100 93.100 39.950 ;
        RECT 19.150 6.700 93.100 7.100 ;
        RECT 19.150 6.600 23.500 6.700 ;
        RECT 7.450 -0.635 10.000 -0.630 ;
        RECT -9.210 -0.805 -7.370 -0.635 ;
        RECT -5.770 -0.805 3.890 -0.635 ;
        RECT 5.700 -0.805 10.000 -0.635 ;
        RECT -8.650 -1.565 -8.320 -0.805 ;
        RECT -7.720 -1.955 -7.460 -0.805 ;
        RECT -6.750 -1.580 -6.350 -1.080 ;
        RECT -5.255 -1.305 -4.925 -0.805 ;
        RECT -4.315 -1.305 -3.985 -0.805 ;
        RECT -2.340 -1.185 -1.960 -0.805 ;
        RECT -1.440 -1.185 -1.110 -0.805 ;
        RECT 0.170 -1.185 0.590 -0.805 ;
        RECT 1.260 -1.495 1.590 -0.805 ;
        RECT 2.710 -1.605 2.995 -0.805 ;
        RECT 6.260 -1.565 6.590 -0.805 ;
        RECT 7.190 -0.980 10.000 -0.805 ;
        RECT 7.190 -1.955 7.450 -0.980 ;
        RECT 9.650 -1.430 10.000 -0.980 ;
        RECT -7.850 -5.845 -0.700 -5.830 ;
        RECT -9.060 -6.015 -0.700 -5.845 ;
        RECT -9.750 -6.630 -9.350 -6.130 ;
        RECT -8.935 -7.155 -8.705 -6.015 ;
        RECT -8.035 -6.180 -0.700 -6.015 ;
        RECT -8.035 -7.155 -7.825 -6.180 ;
        RECT -1.050 -6.315 -0.700 -6.180 ;
        RECT -1.050 -6.485 2.170 -6.315 ;
        RECT 3.530 -6.330 5.370 -6.315 ;
        RECT 9.650 -6.330 10.000 -5.880 ;
        RECT 3.530 -6.485 10.000 -6.330 ;
        RECT 0.005 -7.335 0.175 -6.485 ;
        RECT 0.845 -6.995 1.015 -6.485 ;
        RECT 2.700 -7.380 3.100 -6.880 ;
        RECT 4.090 -7.245 4.420 -6.485 ;
        RECT 5.020 -6.680 10.000 -6.485 ;
        RECT 5.020 -7.635 5.280 -6.680 ;
        RECT 9.650 -7.080 10.000 -6.680 ;
        RECT 42.440 -7.125 44.740 -6.955 ;
        RECT 41.800 -7.970 42.100 -7.470 ;
        RECT 42.955 -7.525 43.890 -7.125 ;
        RECT 44.415 -8.450 44.655 -7.805 ;
        RECT 44.415 -8.750 44.800 -8.450 ;
        RECT 44.415 -8.785 44.655 -8.750 ;
        RECT -8.055 -13.725 -7.845 -12.585 ;
        RECT -7.175 -13.725 -6.945 -12.585 ;
        RECT -6.350 -13.330 -5.950 -12.830 ;
        RECT -4.835 -13.725 -4.550 -12.925 ;
        RECT -3.430 -13.725 -3.100 -13.035 ;
        RECT -2.430 -13.725 -2.010 -13.345 ;
        RECT -0.730 -13.725 -0.400 -13.345 ;
        RECT 0.120 -13.725 0.500 -13.345 ;
        RECT 2.145 -13.725 2.475 -13.225 ;
        RECT 3.085 -13.725 3.415 -13.225 ;
        RECT 5.950 -13.725 6.210 -12.575 ;
        RECT 6.810 -13.725 7.140 -12.965 ;
        RECT 9.650 -13.680 10.000 -13.230 ;
        RECT 7.650 -13.725 10.000 -13.680 ;
        RECT -8.200 -13.895 -6.820 -13.725 ;
        RECT -5.730 -13.895 3.930 -13.725 ;
        RECT 5.860 -13.895 10.000 -13.725 ;
        RECT 7.650 -14.030 10.000 -13.895 ;
        RECT -7.400 -19.655 -7.000 -19.500 ;
        RECT -7.410 -19.825 -3.730 -19.655 ;
        RECT -3.310 -19.825 0.370 -19.655 ;
        RECT 0.790 -19.825 4.470 -19.655 ;
        RECT 5.190 -19.825 8.870 -19.655 ;
        RECT 9.290 -19.825 12.970 -19.655 ;
        RECT 13.390 -19.825 17.070 -19.655 ;
        RECT -6.755 -20.285 -6.485 -19.825 ;
        RECT -4.695 -20.285 -4.370 -19.825 ;
        RECT -2.655 -20.285 -2.385 -19.825 ;
        RECT -0.595 -20.285 -0.270 -19.825 ;
        RECT 1.445 -20.285 1.715 -19.825 ;
        RECT 3.505 -20.285 3.830 -19.825 ;
        RECT 4.700 -20.650 5.100 -20.150 ;
        RECT 5.845 -20.285 6.115 -19.825 ;
        RECT 7.905 -20.285 8.230 -19.825 ;
        RECT 9.945 -20.285 10.215 -19.825 ;
        RECT 12.005 -20.285 12.330 -19.825 ;
        RECT 14.045 -20.285 14.315 -19.825 ;
        RECT 16.105 -20.285 16.430 -19.825 ;
        RECT 60.040 -20.400 61.880 -20.355 ;
        RECT 65.800 -20.400 66.250 -19.000 ;
        RECT 60.040 -20.525 66.250 -20.400 ;
        RECT 60.600 -21.285 60.930 -20.525 ;
        RECT 61.530 -20.750 66.250 -20.525 ;
        RECT 61.530 -21.675 61.790 -20.750 ;
        RECT 62.150 -21.600 62.450 -20.750 ;
        RECT -5.950 -23.655 -3.200 -23.500 ;
        RECT -7.410 -23.700 3.750 -23.655 ;
        RECT -7.410 -23.825 -5.570 -23.700 ;
        RECT -6.850 -24.585 -6.520 -23.825 ;
        RECT -5.920 -24.975 -5.660 -23.825 ;
        RECT -5.150 -24.650 -4.750 -23.700 ;
        RECT -3.610 -23.825 3.750 -23.700 ;
        RECT 5.640 -23.825 7.020 -23.655 ;
        RECT 8.290 -23.825 9.670 -23.655 ;
        RECT -3.095 -24.325 -2.765 -23.825 ;
        RECT -2.170 -24.285 -1.905 -23.825 ;
        RECT 0.000 -24.625 0.170 -23.825 ;
        RECT 1.880 -24.325 2.195 -23.825 ;
        RECT 2.935 -24.835 3.105 -23.825 ;
        RECT 5.725 -24.965 6.005 -23.825 ;
        RECT 6.675 -24.965 6.935 -23.825 ;
        RECT 8.415 -24.965 8.645 -23.825 ;
        RECT 9.315 -24.965 9.525 -23.825 ;
        RECT 37.600 -24.550 44.250 -24.150 ;
        RECT 37.600 -26.550 38.000 -24.550 ;
        RECT 38.300 -27.850 38.700 -24.550 ;
        RECT 41.350 -26.500 41.750 -24.550 ;
        RECT 42.050 -27.850 42.450 -26.050 ;
        RECT 43.850 -27.850 44.250 -24.550 ;
        RECT 65.850 -25.150 66.250 -20.750 ;
        RECT 79.700 -24.255 81.050 -24.100 ;
        RECT 67.790 -24.425 70.090 -24.255 ;
        RECT 72.390 -24.425 81.050 -24.255 ;
        RECT 67.920 -25.565 68.185 -24.425 ;
        RECT 68.855 -25.225 69.025 -24.425 ;
        RECT 69.695 -24.885 69.905 -24.425 ;
        RECT 72.905 -24.925 73.235 -24.425 ;
        RECT 73.830 -24.885 74.095 -24.425 ;
        RECT 76.000 -25.225 76.170 -24.425 ;
        RECT 77.880 -24.925 78.195 -24.425 ;
        RECT 78.935 -25.435 79.105 -24.425 ;
        RECT 79.700 -24.450 81.050 -24.425 ;
        RECT 80.650 -28.200 81.050 -24.450 ;
        RECT 61.800 -28.900 62.300 -28.300 ;
        RECT 68.350 -28.455 70.000 -28.300 ;
        RECT 65.590 -28.625 70.000 -28.455 ;
        RECT 70.990 -28.625 80.650 -28.455 ;
        RECT 61.800 -29.400 62.900 -28.900 ;
        RECT 64.850 -29.400 65.250 -28.900 ;
        RECT 7.450 -32.285 10.000 -32.280 ;
        RECT -9.210 -32.455 -7.370 -32.285 ;
        RECT -5.770 -32.455 3.890 -32.285 ;
        RECT 5.700 -32.455 10.000 -32.285 ;
        RECT -8.650 -33.215 -8.320 -32.455 ;
        RECT -7.720 -33.605 -7.460 -32.455 ;
        RECT -6.750 -33.230 -6.350 -32.730 ;
        RECT -5.255 -32.955 -4.925 -32.455 ;
        RECT -4.315 -32.955 -3.985 -32.455 ;
        RECT -2.340 -32.835 -1.960 -32.455 ;
        RECT -1.440 -32.835 -1.110 -32.455 ;
        RECT 0.170 -32.835 0.590 -32.455 ;
        RECT 1.260 -33.145 1.590 -32.455 ;
        RECT 2.710 -33.255 2.995 -32.455 ;
        RECT 6.260 -33.215 6.590 -32.455 ;
        RECT 7.190 -32.630 10.000 -32.455 ;
        RECT 7.190 -33.605 7.450 -32.630 ;
        RECT 9.650 -33.080 10.000 -32.630 ;
        RECT 33.875 -35.850 34.045 -35.290 ;
        RECT 33.115 -36.180 34.045 -35.850 ;
        RECT 33.875 -36.780 34.045 -36.180 ;
        RECT 32.725 -37.040 34.045 -36.780 ;
        RECT 33.875 -37.130 34.045 -37.040 ;
        RECT 61.800 -36.350 62.300 -29.400 ;
        RECT 66.185 -29.425 66.425 -28.625 ;
        RECT 66.945 -29.425 67.275 -28.625 ;
        RECT 67.785 -29.775 68.115 -28.625 ;
        RECT 68.350 -28.750 70.000 -28.625 ;
        RECT 71.505 -29.125 71.835 -28.625 ;
        RECT 72.430 -29.085 72.695 -28.625 ;
        RECT 74.600 -29.425 74.770 -28.625 ;
        RECT 76.480 -29.125 76.795 -28.625 ;
        RECT 77.540 -29.635 77.710 -28.625 ;
        RECT 78.380 -29.540 78.555 -28.625 ;
        RECT 79.415 -29.765 79.630 -28.625 ;
        RECT 80.305 -29.765 80.555 -28.625 ;
        RECT 81.000 -29.750 81.500 -29.350 ;
        RECT 79.700 -35.955 81.050 -35.800 ;
        RECT 67.790 -36.125 70.090 -35.955 ;
        RECT 72.390 -36.125 81.050 -35.955 ;
        RECT 61.800 -36.850 62.900 -36.350 ;
        RECT 65.850 -36.850 66.250 -36.350 ;
        RECT -7.850 -37.495 -0.700 -37.480 ;
        RECT -9.060 -37.665 -0.700 -37.495 ;
        RECT -9.750 -38.280 -9.350 -37.780 ;
        RECT -8.935 -38.805 -8.705 -37.665 ;
        RECT -8.035 -37.830 -0.700 -37.665 ;
        RECT -8.035 -38.805 -7.825 -37.830 ;
        RECT -1.050 -37.965 -0.700 -37.830 ;
        RECT -1.050 -38.135 2.170 -37.965 ;
        RECT 3.530 -37.980 5.370 -37.965 ;
        RECT 9.650 -37.980 10.000 -37.530 ;
        RECT 32.900 -37.750 33.400 -37.350 ;
        RECT 61.800 -37.450 62.300 -36.850 ;
        RECT 67.920 -37.265 68.185 -36.125 ;
        RECT 68.855 -36.925 69.025 -36.125 ;
        RECT 69.695 -36.585 69.905 -36.125 ;
        RECT 72.905 -36.625 73.235 -36.125 ;
        RECT 73.830 -36.585 74.095 -36.125 ;
        RECT 76.000 -36.925 76.170 -36.125 ;
        RECT 77.880 -36.625 78.195 -36.125 ;
        RECT 78.935 -37.135 79.105 -36.125 ;
        RECT 79.700 -36.150 81.050 -36.125 ;
        RECT 3.530 -38.135 10.000 -37.980 ;
        RECT 0.005 -38.985 0.175 -38.135 ;
        RECT 0.845 -38.645 1.015 -38.135 ;
        RECT 2.700 -39.030 3.100 -38.530 ;
        RECT 4.090 -38.895 4.420 -38.135 ;
        RECT 5.020 -38.330 10.000 -38.135 ;
        RECT 5.020 -39.285 5.280 -38.330 ;
        RECT 9.650 -38.730 10.000 -38.330 ;
        RECT 33.875 -38.715 34.045 -38.590 ;
        RECT 32.735 -38.945 34.045 -38.715 ;
        RECT 33.875 -39.615 34.045 -38.945 ;
        RECT 32.735 -39.825 34.045 -39.615 ;
        RECT 33.875 -39.970 34.045 -39.825 ;
        RECT 80.650 -39.900 81.050 -36.150 ;
        RECT 68.350 -40.155 70.000 -40.000 ;
        RECT 65.590 -40.325 70.000 -40.155 ;
        RECT 70.990 -40.325 80.650 -40.155 ;
        RECT 64.850 -41.100 65.250 -40.600 ;
        RECT 66.185 -41.125 66.425 -40.325 ;
        RECT 66.945 -41.125 67.275 -40.325 ;
        RECT 67.785 -41.475 68.115 -40.325 ;
        RECT 68.350 -40.450 70.000 -40.325 ;
        RECT 71.505 -40.825 71.835 -40.325 ;
        RECT 72.430 -40.785 72.695 -40.325 ;
        RECT 74.600 -41.125 74.770 -40.325 ;
        RECT 76.480 -40.825 76.795 -40.325 ;
        RECT 77.540 -41.335 77.710 -40.325 ;
        RECT 78.380 -41.240 78.555 -40.325 ;
        RECT 79.415 -41.465 79.630 -40.325 ;
        RECT 80.305 -41.465 80.555 -40.325 ;
        RECT 81.000 -41.450 81.500 -41.050 ;
        RECT -8.055 -45.375 -7.845 -44.235 ;
        RECT -7.175 -45.375 -6.945 -44.235 ;
        RECT -6.350 -44.980 -5.950 -44.480 ;
        RECT -4.835 -45.375 -4.550 -44.575 ;
        RECT -3.430 -45.375 -3.100 -44.685 ;
        RECT -2.430 -45.375 -2.010 -44.995 ;
        RECT -0.730 -45.375 -0.400 -44.995 ;
        RECT 0.120 -45.375 0.500 -44.995 ;
        RECT 2.145 -45.375 2.475 -44.875 ;
        RECT 3.085 -45.375 3.415 -44.875 ;
        RECT 5.950 -45.375 6.210 -44.225 ;
        RECT 6.810 -45.375 7.140 -44.615 ;
        RECT 9.650 -45.330 10.000 -44.880 ;
        RECT 7.650 -45.375 10.000 -45.330 ;
        RECT -8.200 -45.400 -6.820 -45.375 ;
        RECT -15.300 -45.545 -6.820 -45.400 ;
        RECT -5.730 -45.545 3.930 -45.375 ;
        RECT 5.860 -45.545 10.000 -45.375 ;
        RECT -15.300 -46.400 -7.700 -45.545 ;
        RECT 7.650 -45.680 10.000 -45.545 ;
      LAYER met1 ;
        RECT -1.450 39.950 0.550 40.350 ;
        RECT 15.100 39.950 17.100 40.350 ;
        RECT 55.200 39.950 57.200 40.350 ;
        RECT 79.350 39.950 81.350 40.350 ;
        RECT -6.900 38.600 -6.500 39.100 ;
        RECT 2.600 38.600 3.000 39.100 ;
        RECT 8.050 38.600 8.450 39.100 ;
        RECT 13.500 38.600 13.900 39.100 ;
        RECT 23.100 38.600 23.500 39.100 ;
        RECT 32.600 38.600 33.000 39.100 ;
        RECT 38.050 38.600 38.450 39.100 ;
        RECT 43.500 38.600 43.900 39.100 ;
        RECT 53.100 38.600 53.500 39.100 ;
        RECT 62.600 38.600 63.000 39.100 ;
        RECT 68.050 38.600 68.450 39.100 ;
        RECT 73.500 38.600 73.900 39.100 ;
        RECT 15.450 22.050 19.650 22.550 ;
        RECT 15.550 21.350 16.050 22.050 ;
        RECT 15.540 20.870 17.840 21.350 ;
        RECT 18.100 20.250 18.500 22.050 ;
        RECT 17.350 19.850 17.950 20.150 ;
        RECT 19.150 19.850 19.650 22.050 ;
        RECT 17.350 19.550 19.650 19.850 ;
        RECT 31.900 7.950 32.300 8.450 ;
        RECT 37.350 7.950 37.750 8.450 ;
        RECT 42.800 7.950 43.200 8.450 ;
        RECT 52.300 7.950 52.700 8.450 ;
        RECT 61.900 7.950 62.300 8.450 ;
        RECT 67.350 7.950 67.750 8.450 ;
        RECT 72.800 7.950 73.200 8.450 ;
        RECT 82.300 7.950 82.700 8.450 ;
        RECT -7.400 -0.480 -5.400 5.550 ;
        RECT -1.600 -0.480 0.400 5.550 ;
        RECT 4.450 -0.480 6.450 5.550 ;
        RECT -9.210 -0.960 7.540 -0.480 ;
        RECT -7.400 -0.980 -5.700 -0.960 ;
        RECT 3.850 -0.980 5.700 -0.960 ;
        RECT 9.200 -0.980 10.000 -0.630 ;
        RECT -6.750 -1.580 -6.350 -0.980 ;
        RECT -9.750 -5.690 -9.000 -5.680 ;
        RECT -9.750 -6.170 -7.680 -5.690 ;
        RECT 2.150 -6.160 3.550 -6.130 ;
        RECT -9.750 -6.180 -9.000 -6.170 ;
        RECT -9.750 -6.630 -9.350 -6.180 ;
        RECT -1.050 -6.630 5.370 -6.160 ;
        RECT -1.050 -6.640 2.170 -6.630 ;
        RECT 2.700 -7.380 3.100 -6.630 ;
        RECT 3.530 -6.640 5.370 -6.630 ;
        RECT -8.200 -13.580 -6.820 -13.570 ;
        RECT -6.350 -13.580 -5.950 -12.830 ;
        RECT -5.730 -13.580 3.930 -13.570 ;
        RECT 5.860 -13.580 7.700 -13.570 ;
        RECT -8.200 -14.030 7.700 -13.580 ;
        RECT 9.650 -13.680 10.000 -0.980 ;
        RECT 37.100 -7.250 45.600 -6.800 ;
        RECT 41.800 -7.970 42.100 -7.250 ;
        RECT 42.440 -7.280 44.740 -7.250 ;
        RECT 45.250 -8.450 45.600 -7.250 ;
        RECT 44.400 -8.800 45.600 -8.450 ;
        RECT 9.250 -14.030 10.000 -13.680 ;
        RECT -8.200 -14.050 -6.820 -14.030 ;
        RECT -5.730 -14.050 3.930 -14.030 ;
        RECT 5.860 -14.050 7.700 -14.030 ;
        RECT 65.800 -19.000 66.250 -17.700 ;
        RECT 65.200 -19.450 66.250 -19.000 ;
        RECT -11.600 -19.980 17.070 -19.500 ;
        RECT -11.600 -20.000 -7.300 -19.980 ;
        RECT -3.750 -20.000 -3.250 -19.980 ;
        RECT 0.350 -20.000 0.850 -19.980 ;
        RECT 4.450 -20.000 5.200 -19.980 ;
        RECT 8.850 -20.000 9.300 -19.980 ;
        RECT 12.950 -20.000 13.400 -19.980 ;
        RECT -11.600 -23.500 -9.600 -20.000 ;
        RECT 4.700 -20.650 5.100 -20.000 ;
        RECT 60.040 -20.680 61.880 -20.200 ;
        RECT 62.150 -21.600 62.450 -21.100 ;
        RECT -11.600 -23.980 -5.570 -23.500 ;
        RECT -3.610 -23.980 9.670 -23.500 ;
        RECT -11.600 -24.000 -7.300 -23.980 ;
        RECT 3.750 -24.000 5.650 -23.980 ;
        RECT 7.000 -24.000 8.300 -23.980 ;
        RECT -5.150 -24.650 -4.750 -24.150 ;
        RECT 33.700 -24.550 38.700 -24.150 ;
        RECT -9.210 -32.610 7.540 -32.130 ;
        RECT -7.400 -32.630 -5.700 -32.610 ;
        RECT 3.850 -32.630 5.700 -32.610 ;
        RECT 9.200 -32.630 10.000 -32.280 ;
        RECT -6.750 -33.230 -6.350 -32.630 ;
        RECT -9.750 -37.340 -9.000 -37.330 ;
        RECT -9.750 -37.820 -7.680 -37.340 ;
        RECT 2.150 -37.810 3.550 -37.780 ;
        RECT -9.750 -37.830 -9.000 -37.820 ;
        RECT -9.750 -38.280 -9.350 -37.830 ;
        RECT -1.050 -38.280 5.370 -37.810 ;
        RECT -1.050 -38.290 2.170 -38.280 ;
        RECT 2.700 -39.030 3.100 -38.280 ;
        RECT 3.530 -38.290 5.370 -38.280 ;
        RECT -8.200 -45.230 -6.820 -45.220 ;
        RECT -6.350 -45.230 -5.950 -44.480 ;
        RECT -5.730 -45.230 3.930 -45.220 ;
        RECT 5.860 -45.230 7.700 -45.220 ;
        RECT -15.300 -46.400 -12.900 -45.400 ;
        RECT -8.200 -45.680 7.700 -45.230 ;
        RECT 9.650 -45.330 10.000 -32.630 ;
        RECT 33.700 -35.300 34.200 -24.550 ;
        RECT 67.790 -24.580 79.750 -24.100 ;
        RECT 70.050 -24.600 72.500 -24.580 ;
        RECT 61.800 -25.150 66.250 -24.650 ;
        RECT 37.600 -26.550 38.000 -26.050 ;
        RECT 41.350 -26.500 41.750 -26.000 ;
        RECT 42.050 -26.200 42.450 -26.050 ;
        RECT 43.850 -26.200 44.250 -26.050 ;
        RECT 42.050 -26.700 44.250 -26.200 ;
        RECT 42.050 -26.850 42.450 -26.700 ;
        RECT 43.850 -26.850 44.250 -26.700 ;
        RECT 61.800 -28.900 62.300 -25.150 ;
        RECT 80.650 -28.300 81.050 -27.800 ;
        RECT 64.850 -28.750 68.350 -28.300 ;
        RECT 69.500 -28.750 81.050 -28.300 ;
        RECT 64.850 -28.900 65.250 -28.750 ;
        RECT 65.590 -28.780 68.350 -28.750 ;
        RECT 70.990 -28.780 81.050 -28.750 ;
        RECT 80.650 -28.800 81.050 -28.780 ;
        RECT 61.800 -29.400 65.250 -28.900 ;
        RECT 81.000 -29.750 81.500 -29.350 ;
        RECT 33.720 -37.100 34.200 -35.300 ;
        RECT 67.790 -36.280 79.750 -35.800 ;
        RECT 70.050 -36.300 72.500 -36.280 ;
        RECT 33.700 -37.350 34.200 -37.100 ;
        RECT 32.900 -37.750 34.200 -37.350 ;
        RECT 33.700 -38.600 34.200 -37.750 ;
        RECT 33.720 -39.970 34.200 -38.600 ;
        RECT 61.800 -36.850 66.250 -36.350 ;
        RECT 61.800 -40.600 62.300 -36.850 ;
        RECT 80.650 -40.000 81.050 -39.500 ;
        RECT 64.850 -40.450 68.350 -40.000 ;
        RECT 69.500 -40.450 81.050 -40.000 ;
        RECT 64.850 -40.600 65.250 -40.450 ;
        RECT 65.590 -40.480 68.350 -40.450 ;
        RECT 70.990 -40.480 81.050 -40.450 ;
        RECT 80.650 -40.500 81.050 -40.480 ;
        RECT 61.250 -41.100 65.250 -40.600 ;
        RECT 81.000 -41.450 81.500 -41.050 ;
        RECT 9.250 -45.680 10.000 -45.330 ;
        RECT -8.200 -45.700 -6.200 -45.680 ;
        RECT -5.730 -45.700 4.900 -45.680 ;
        RECT 5.860 -45.700 7.700 -45.680 ;
        RECT 2.900 -46.250 4.900 -45.700 ;
        RECT -15.300 -47.950 -13.300 -46.400 ;
      LAYER met2 ;
        RECT -1.450 39.950 0.550 41.050 ;
        RECT 15.100 39.950 17.100 41.050 ;
        RECT 55.200 39.950 57.200 41.100 ;
        RECT 79.350 39.950 81.350 41.050 ;
        RECT -7.400 3.550 -5.400 5.550 ;
        RECT -1.600 3.550 0.400 5.550 ;
        RECT 4.450 3.550 6.450 5.550 ;
        RECT 37.100 -19.000 37.600 -6.800 ;
        RECT 65.800 -19.000 67.100 -17.700 ;
        RECT 37.100 -19.450 67.100 -19.000 ;
        RECT -11.600 -22.950 -9.600 -20.950 ;
        RECT 37.100 -24.550 37.600 -19.450 ;
        RECT 65.800 -19.700 67.100 -19.450 ;
        RECT 61.250 -41.600 63.250 -40.600 ;
        RECT 2.900 -46.800 4.900 -45.700 ;
        RECT -15.300 -47.950 -13.300 -46.850 ;
      LAYER met3 ;
        RECT -31.620 56.780 114.600 59.500 ;
        RECT -1.450 40.350 0.550 41.050 ;
        RECT 15.100 40.350 17.100 41.850 ;
        RECT 55.200 40.350 57.200 41.850 ;
        RECT 79.350 40.350 81.350 41.750 ;
        RECT -31.450 3.550 6.450 5.550 ;
        RECT 65.800 -19.700 114.600 -17.700 ;
        RECT -31.450 -22.950 -9.600 -20.950 ;
        RECT 61.250 -42.200 63.250 -41.100 ;
        RECT -15.300 -48.600 -13.300 -47.300 ;
        RECT 2.900 -47.400 4.900 -46.200 ;
        RECT -31.620 -70.380 114.600 -67.660 ;
      LAYER met4 ;
        RECT -31.620 -70.380 -28.900 59.500 ;
        RECT -1.500 58.950 0.500 59.500 ;
        RECT -1.500 56.700 0.550 58.950 ;
        RECT -1.500 41.300 0.500 56.700 ;
        RECT -1.500 41.200 0.550 41.300 ;
        RECT -1.450 39.950 0.550 41.200 ;
        RECT 15.100 39.950 17.100 58.950 ;
        RECT 55.200 39.950 57.200 58.950 ;
        RECT 79.350 39.950 81.350 58.950 ;
        RECT 111.880 56.700 114.600 59.500 ;
        RECT 111.900 -17.700 114.600 56.700 ;
        RECT 111.880 -19.700 114.600 -17.700 ;
        RECT -15.300 -48.500 -13.300 -46.850 ;
        RECT -15.300 -70.400 -13.200 -48.500 ;
        RECT 2.900 -70.350 4.900 -45.700 ;
        RECT 61.250 -70.350 63.250 -40.600 ;
        RECT 111.900 -67.600 114.600 -19.700 ;
        RECT 111.880 -70.380 114.600 -67.600 ;
    END
  END VDDA
  PIN GND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -7.100 28.600 82.900 33.400 ;
        RECT 16.030 19.400 17.835 19.405 ;
        RECT 16.030 19.175 18.750 19.400 ;
        RECT 15.545 18.500 18.750 19.175 ;
        RECT 15.545 18.495 17.835 18.500 ;
        RECT 15.690 18.305 15.860 18.495 ;
        RECT 22.900 13.650 82.900 18.450 ;
        RECT 34.400 -1.150 36.700 -1.050 ;
        RECT 36.900 -1.150 47.600 -1.050 ;
        RECT 47.800 -1.150 52.300 -1.050 ;
        RECT 52.500 -1.150 63.200 -1.050 ;
        RECT 63.400 -1.150 67.900 -1.050 ;
        RECT 68.100 -1.150 78.800 -1.050 ;
        RECT 79.000 -1.150 81.200 -1.050 ;
        RECT -8.720 -2.630 -7.375 -2.425 ;
        RECT -10.000 -2.655 -9.150 -2.630 ;
        RECT -8.720 -2.655 -5.750 -2.630 ;
        RECT -4.405 -2.655 -3.485 -2.435 ;
        RECT 2.595 -2.535 3.515 -2.425 ;
        RECT 1.180 -2.630 3.515 -2.535 ;
        RECT 1.180 -2.655 5.750 -2.630 ;
        RECT 6.190 -2.655 7.535 -2.425 ;
        RECT -10.000 -3.330 7.535 -2.655 ;
        RECT -9.205 -3.335 -7.375 -3.330 ;
        RECT -5.765 -3.335 3.515 -3.330 ;
        RECT 5.705 -3.335 7.535 -3.330 ;
        RECT -9.065 -3.525 -8.895 -3.335 ;
        RECT -5.625 -3.525 -5.455 -3.335 ;
        RECT 5.845 -3.525 6.015 -3.335 ;
        RECT 34.400 -3.850 81.200 -1.150 ;
        RECT -9.950 -7.635 -9.000 -7.630 ;
        RECT -9.950 -8.530 -7.695 -7.635 ;
        RECT -9.045 -8.545 -7.695 -8.530 ;
        RECT -1.005 -8.330 2.165 -8.105 ;
        RECT -1.005 -8.335 3.550 -8.330 ;
        RECT 4.020 -8.335 5.365 -8.105 ;
        RECT -8.915 -8.735 -8.745 -8.545 ;
        RECT -1.005 -9.015 5.365 -8.335 ;
        RECT 42.930 -8.975 44.735 -8.745 ;
        RECT 42.445 -8.980 44.735 -8.975 ;
        RECT -0.905 -9.205 -0.735 -9.015 ;
        RECT 2.150 -9.030 3.550 -9.015 ;
        RECT 3.675 -9.205 3.845 -9.015 ;
        RECT 41.780 -9.655 44.735 -8.980 ;
        RECT 41.780 -9.660 42.450 -9.655 ;
        RECT 42.590 -9.845 42.760 -9.655 ;
        RECT -7.135 -11.195 -6.965 -11.005 ;
        RECT -6.850 -11.195 -5.350 -11.180 ;
        RECT 3.615 -11.195 3.785 -11.005 ;
        RECT 3.900 -11.195 5.900 -11.180 ;
        RECT 7.385 -11.195 7.555 -11.005 ;
        RECT -8.185 -11.875 7.695 -11.195 ;
        RECT -8.185 -11.995 -3.020 -11.875 ;
        RECT -8.185 -12.105 -4.435 -11.995 ;
        RECT 1.645 -12.095 2.565 -11.875 ;
        RECT 3.900 -11.880 7.210 -11.875 ;
        RECT 5.865 -12.105 7.210 -11.880 ;
        RECT 48.850 -11.950 80.050 -9.250 ;
        RECT 48.850 -12.050 51.050 -11.950 ;
        RECT 51.250 -12.050 61.950 -11.950 ;
        RECT 62.150 -12.050 66.650 -11.950 ;
        RECT 66.850 -12.050 77.550 -11.950 ;
        RECT 77.750 -12.050 80.050 -11.950 ;
        RECT -6.850 -12.130 -5.350 -12.105 ;
        RECT -7.600 -22.400 17.300 -21.400 ;
        RECT 60.530 -22.150 61.875 -22.145 ;
        RECT 60.530 -22.375 62.700 -22.150 ;
        RECT -7.265 -22.545 -7.095 -22.400 ;
        RECT -3.165 -22.545 -2.995 -22.400 ;
        RECT 0.935 -22.545 1.105 -22.400 ;
        RECT 5.335 -22.545 5.505 -22.400 ;
        RECT 9.435 -22.545 9.605 -22.400 ;
        RECT 13.535 -22.545 13.705 -22.400 ;
        RECT 60.045 -23.050 62.700 -22.375 ;
        RECT 60.045 -23.055 61.875 -23.050 ;
        RECT 60.185 -23.245 60.355 -23.055 ;
        RECT -7.600 -26.400 9.900 -25.400 ;
        RECT 65.550 -26.045 67.900 -26.000 ;
        RECT 65.550 -26.250 70.035 -26.045 ;
        RECT 65.550 -26.275 72.450 -26.250 ;
        RECT 75.910 -26.275 76.820 -26.055 ;
        RECT 78.355 -26.275 79.705 -26.045 ;
        RECT -7.265 -26.545 -7.095 -26.400 ;
        RECT -3.465 -26.545 -3.295 -26.400 ;
        RECT 5.780 -26.545 5.950 -26.400 ;
        RECT 8.435 -26.545 8.605 -26.400 ;
        RECT 65.550 -26.955 79.705 -26.275 ;
        RECT 65.550 -27.000 67.900 -26.955 ;
        RECT 67.935 -27.145 68.105 -26.955 ;
        RECT 70.000 -27.000 72.450 -26.955 ;
        RECT 72.535 -27.145 72.705 -26.955 ;
        RECT 65.595 -30.250 68.205 -30.245 ;
        RECT 64.550 -30.450 68.205 -30.250 ;
        RECT 64.550 -30.475 71.050 -30.450 ;
        RECT 74.510 -30.475 75.420 -30.255 ;
        RECT 76.960 -30.475 80.645 -30.245 ;
        RECT 64.550 -31.155 80.645 -30.475 ;
        RECT 64.550 -31.500 65.650 -31.155 ;
        RECT 65.740 -31.345 65.910 -31.155 ;
        RECT 68.200 -31.200 71.050 -31.155 ;
        RECT 71.135 -31.345 71.305 -31.155 ;
        RECT -8.720 -34.280 -7.375 -34.075 ;
        RECT -10.000 -34.305 -9.150 -34.280 ;
        RECT -8.720 -34.305 -5.750 -34.280 ;
        RECT -4.405 -34.305 -3.485 -34.085 ;
        RECT 2.595 -34.185 3.515 -34.075 ;
        RECT 1.180 -34.280 3.515 -34.185 ;
        RECT 1.180 -34.305 5.750 -34.280 ;
        RECT 6.190 -34.305 7.535 -34.075 ;
        RECT -10.000 -34.980 7.535 -34.305 ;
        RECT -9.205 -34.985 -7.375 -34.980 ;
        RECT -5.765 -34.985 3.515 -34.980 ;
        RECT 5.705 -34.985 7.535 -34.980 ;
        RECT -9.065 -35.175 -8.895 -34.985 ;
        RECT -5.625 -35.175 -5.455 -34.985 ;
        RECT 5.845 -35.175 6.015 -34.985 ;
        RECT 31.345 -35.435 32.025 -35.295 ;
        RECT 31.155 -35.605 32.025 -35.435 ;
        RECT 31.345 -35.780 32.025 -35.605 ;
        RECT 42.550 -35.650 45.850 -32.850 ;
        RECT 47.100 -35.650 50.400 -32.850 ;
        RECT 31.345 -37.125 32.255 -35.780 ;
        RECT 31.350 -38.605 32.250 -37.125 ;
        RECT 65.550 -37.745 67.900 -37.700 ;
        RECT 65.550 -37.950 70.035 -37.745 ;
        RECT 65.550 -37.975 72.450 -37.950 ;
        RECT 75.910 -37.975 76.820 -37.755 ;
        RECT 78.355 -37.975 79.705 -37.745 ;
        RECT 31.345 -38.735 32.255 -38.605 ;
        RECT 65.550 -38.655 79.705 -37.975 ;
        RECT 65.550 -38.700 67.900 -38.655 ;
        RECT 31.155 -38.905 32.255 -38.735 ;
        RECT 67.935 -38.845 68.105 -38.655 ;
        RECT 70.000 -38.700 72.450 -38.655 ;
        RECT 72.535 -38.845 72.705 -38.655 ;
        RECT -9.950 -39.285 -9.000 -39.280 ;
        RECT -9.950 -40.180 -7.695 -39.285 ;
        RECT -9.045 -40.195 -7.695 -40.180 ;
        RECT -1.005 -39.980 2.165 -39.755 ;
        RECT -1.005 -39.985 3.550 -39.980 ;
        RECT 4.020 -39.985 5.365 -39.755 ;
        RECT 31.345 -39.955 32.255 -38.905 ;
        RECT -8.915 -40.385 -8.745 -40.195 ;
        RECT -1.005 -40.665 5.365 -39.985 ;
        RECT -0.905 -40.855 -0.735 -40.665 ;
        RECT 2.150 -40.680 3.550 -40.665 ;
        RECT 3.675 -40.855 3.845 -40.665 ;
        RECT -7.135 -42.845 -6.965 -42.655 ;
        RECT -6.850 -42.845 -5.350 -42.830 ;
        RECT 3.615 -42.845 3.785 -42.655 ;
        RECT 3.900 -42.845 5.900 -42.830 ;
        RECT 7.385 -42.845 7.555 -42.655 ;
        RECT -8.185 -43.525 7.695 -42.845 ;
        RECT -8.185 -43.645 -3.020 -43.525 ;
        RECT -8.185 -43.755 -4.435 -43.645 ;
        RECT 1.645 -43.745 2.565 -43.525 ;
        RECT 3.900 -43.530 7.210 -43.525 ;
        RECT 5.865 -43.755 7.210 -43.530 ;
        RECT 40.000 -43.650 54.380 -41.640 ;
        RECT 65.595 -41.950 68.205 -41.945 ;
        RECT 64.550 -42.150 68.205 -41.950 ;
        RECT 64.550 -42.175 71.050 -42.150 ;
        RECT 74.510 -42.175 75.420 -41.955 ;
        RECT 76.960 -42.175 80.645 -41.945 ;
        RECT 64.550 -42.855 80.645 -42.175 ;
        RECT 64.550 -43.200 65.650 -42.855 ;
        RECT 65.740 -43.045 65.910 -42.855 ;
        RECT 68.200 -42.900 71.050 -42.855 ;
        RECT 71.135 -43.045 71.305 -42.855 ;
        RECT -6.850 -43.780 -5.350 -43.755 ;
      LAYER li1 ;
        RECT -6.900 28.950 -6.500 29.450 ;
        RECT 2.600 28.950 3.000 29.450 ;
        RECT 8.050 28.950 8.450 29.450 ;
        RECT 13.500 28.950 13.900 29.450 ;
        RECT 23.100 28.950 23.500 29.450 ;
        RECT 32.600 28.950 33.000 29.450 ;
        RECT 38.050 28.950 38.450 29.450 ;
        RECT 43.500 28.950 43.900 29.450 ;
        RECT 53.100 28.950 53.500 29.450 ;
        RECT 62.600 28.950 63.000 29.450 ;
        RECT 68.050 28.950 68.450 29.450 ;
        RECT 73.500 28.950 73.900 29.450 ;
        RECT 31.000 23.050 31.170 23.130 ;
        RECT 29.185 22.730 31.170 23.050 ;
        RECT 31.000 22.650 31.170 22.730 ;
        RECT 16.055 18.475 16.990 18.875 ;
        RECT 18.100 18.750 18.500 19.250 ;
        RECT 15.540 18.305 17.840 18.475 ;
        RECT 31.900 17.600 32.300 18.100 ;
        RECT 37.350 17.600 37.750 18.100 ;
        RECT 42.800 17.600 43.200 18.100 ;
        RECT 52.300 17.600 52.700 18.100 ;
        RECT 61.900 17.600 62.300 18.100 ;
        RECT 67.350 17.600 67.750 18.100 ;
        RECT 72.800 17.600 73.200 18.100 ;
        RECT 82.300 17.600 82.700 18.100 ;
        RECT -9.800 -3.180 -9.400 -2.680 ;
        RECT -8.650 -3.355 -8.320 -2.975 ;
        RECT -7.720 -3.180 -7.460 -2.515 ;
        RECT -7.720 -3.355 -5.750 -3.180 ;
        RECT -5.255 -3.355 -4.925 -2.975 ;
        RECT -4.315 -3.355 -3.985 -2.975 ;
        RECT -2.160 -3.355 -1.750 -2.915 ;
        RECT -1.010 -3.355 -0.690 -2.895 ;
        RECT 0.920 -3.355 1.580 -2.875 ;
        RECT 2.710 -3.355 2.995 -2.895 ;
        RECT 3.850 -3.355 5.700 -3.230 ;
        RECT 6.260 -3.355 6.590 -2.975 ;
        RECT 7.190 -3.355 7.450 -2.515 ;
        RECT -9.210 -3.525 7.540 -3.355 ;
        RECT -7.500 -3.680 -5.750 -3.525 ;
        RECT 3.850 -3.680 5.700 -3.525 ;
        RECT 34.600 -4.350 35.000 -3.000 ;
        RECT 35.300 -4.350 35.700 -1.450 ;
        RECT 38.500 -4.350 38.900 -1.450 ;
        RECT 40.000 -3.000 40.400 -1.450 ;
        RECT 43.100 -3.000 43.500 -1.450 ;
        RECT 39.300 -3.450 40.400 -3.000 ;
        RECT 39.300 -3.500 39.700 -3.450 ;
        RECT 40.000 -4.350 40.400 -3.450 ;
        RECT 42.400 -3.450 43.500 -3.000 ;
        RECT 42.400 -3.500 42.800 -3.450 ;
        RECT 43.100 -4.350 43.500 -3.450 ;
        RECT 45.500 -4.350 45.900 -3.000 ;
        RECT 46.200 -4.350 46.600 -1.450 ;
        RECT 49.400 -4.350 49.800 -1.450 ;
        RECT 50.200 -4.350 50.600 -3.000 ;
        RECT 50.900 -4.350 51.300 -1.450 ;
        RECT 54.100 -4.350 54.500 -1.450 ;
        RECT 55.600 -3.000 56.000 -1.450 ;
        RECT 58.700 -3.000 59.100 -1.450 ;
        RECT 54.900 -3.450 56.000 -3.000 ;
        RECT 54.900 -3.500 55.300 -3.450 ;
        RECT 55.600 -4.350 56.000 -3.450 ;
        RECT 58.000 -3.450 59.100 -3.000 ;
        RECT 58.000 -3.500 58.400 -3.450 ;
        RECT 58.700 -4.350 59.100 -3.450 ;
        RECT 61.100 -4.350 61.500 -3.000 ;
        RECT 61.800 -4.350 62.200 -1.450 ;
        RECT 65.000 -4.350 65.400 -1.450 ;
        RECT 65.800 -4.350 66.200 -3.000 ;
        RECT 66.500 -4.350 66.900 -1.450 ;
        RECT 69.700 -4.350 70.100 -1.450 ;
        RECT 71.200 -3.000 71.600 -1.450 ;
        RECT 74.300 -3.000 74.700 -1.450 ;
        RECT 70.500 -3.450 71.600 -3.000 ;
        RECT 70.500 -3.500 70.900 -3.450 ;
        RECT 71.200 -4.350 71.600 -3.450 ;
        RECT 73.600 -3.450 74.700 -3.000 ;
        RECT 73.600 -3.500 74.000 -3.450 ;
        RECT 74.300 -4.350 74.700 -3.450 ;
        RECT 76.700 -4.350 77.100 -3.000 ;
        RECT 77.400 -4.350 77.800 -1.450 ;
        RECT 80.600 -4.350 81.000 -1.450 ;
        RECT 34.600 -4.750 81.000 -4.350 ;
        RECT -9.750 -8.380 -9.350 -7.880 ;
        RECT -8.935 -8.565 -8.705 -7.745 ;
        RECT -8.035 -8.380 -7.825 -7.745 ;
        RECT -8.035 -8.565 -3.150 -8.380 ;
        RECT -9.060 -8.730 -3.150 -8.565 ;
        RECT -9.060 -8.735 -7.680 -8.730 ;
        RECT -3.500 -8.930 -3.150 -8.730 ;
        RECT -0.915 -8.930 -0.585 -8.645 ;
        RECT -3.500 -9.035 -0.585 -8.930 ;
        RECT -0.075 -9.035 0.255 -8.645 ;
        RECT 1.795 -9.035 2.085 -8.200 ;
        RECT 2.600 -8.880 3.100 -8.480 ;
        RECT 4.090 -9.035 4.420 -8.655 ;
        RECT 5.020 -9.035 5.280 -8.195 ;
        RECT 49.050 -8.350 49.450 -4.750 ;
        RECT 79.450 -8.250 79.850 -4.750 ;
        RECT 79.450 -8.350 93.050 -8.250 ;
        RECT 49.050 -8.750 93.050 -8.350 ;
        RECT -3.500 -9.205 2.170 -9.035 ;
        RECT 3.530 -9.205 5.370 -9.035 ;
        RECT -3.500 -9.280 -0.850 -9.205 ;
        RECT -6.950 -11.005 -5.650 -10.880 ;
        RECT -3.500 -11.005 -3.150 -9.280 ;
        RECT 41.850 -9.600 42.200 -9.050 ;
        RECT 42.955 -9.675 43.890 -9.275 ;
        RECT 42.440 -9.845 44.740 -9.675 ;
        RECT 3.900 -11.005 6.050 -10.980 ;
        RECT 7.350 -11.005 13.700 -10.650 ;
        RECT -8.200 -11.150 13.700 -11.005 ;
        RECT -8.200 -11.175 7.700 -11.150 ;
        RECT -8.055 -11.995 -7.845 -11.175 ;
        RECT -7.175 -11.330 -5.650 -11.175 ;
        RECT -7.175 -11.995 -6.945 -11.330 ;
        RECT -4.835 -11.635 -4.550 -11.175 ;
        RECT -3.420 -11.655 -2.760 -11.175 ;
        RECT -1.150 -11.635 -0.830 -11.175 ;
        RECT -0.090 -11.615 0.320 -11.175 ;
        RECT 2.145 -11.555 2.475 -11.175 ;
        RECT 3.085 -11.555 3.415 -11.175 ;
        RECT 3.900 -11.330 6.210 -11.175 ;
        RECT 5.000 -11.730 5.500 -11.330 ;
        RECT 5.950 -12.015 6.210 -11.330 ;
        RECT 6.810 -11.555 7.140 -11.175 ;
        RECT 49.050 -11.650 49.450 -8.750 ;
        RECT 52.250 -11.650 52.650 -8.750 ;
        RECT 52.950 -10.100 53.350 -8.750 ;
        RECT 55.350 -9.650 55.750 -8.750 ;
        RECT 56.050 -9.650 56.450 -9.600 ;
        RECT 55.350 -10.100 56.450 -9.650 ;
        RECT 58.450 -9.650 58.850 -8.750 ;
        RECT 59.150 -9.650 59.550 -9.600 ;
        RECT 58.450 -10.100 59.550 -9.650 ;
        RECT 55.350 -11.650 55.750 -10.100 ;
        RECT 58.450 -11.650 58.850 -10.100 ;
        RECT 59.950 -11.650 60.350 -8.750 ;
        RECT 63.150 -11.650 63.550 -8.750 ;
        RECT 63.850 -10.100 64.250 -8.750 ;
        RECT 64.650 -11.650 65.050 -8.750 ;
        RECT 67.850 -11.650 68.250 -8.750 ;
        RECT 68.550 -10.100 68.950 -8.750 ;
        RECT 70.950 -9.650 71.350 -8.750 ;
        RECT 71.650 -9.650 72.050 -9.600 ;
        RECT 70.950 -10.100 72.050 -9.650 ;
        RECT 74.050 -9.650 74.450 -8.750 ;
        RECT 74.750 -9.650 75.150 -9.600 ;
        RECT 74.050 -10.100 75.150 -9.650 ;
        RECT 70.950 -11.650 71.350 -10.100 ;
        RECT 74.050 -11.650 74.450 -10.100 ;
        RECT 75.550 -11.650 75.950 -8.750 ;
        RECT 78.750 -11.650 79.150 -8.750 ;
        RECT 79.450 -10.100 79.850 -8.750 ;
        RECT 92.550 -9.350 93.050 -8.750 ;
        RECT -6.755 -22.375 -6.485 -21.915 ;
        RECT -4.695 -22.375 -4.370 -21.915 ;
        RECT -2.655 -22.375 -2.385 -21.915 ;
        RECT -0.595 -22.375 -0.270 -21.915 ;
        RECT 1.445 -22.375 1.715 -21.915 ;
        RECT 3.505 -22.375 3.830 -21.915 ;
        RECT 4.650 -22.210 4.960 -21.710 ;
        RECT 5.845 -22.375 6.115 -21.915 ;
        RECT 7.905 -22.375 8.230 -21.915 ;
        RECT 9.945 -22.375 10.215 -21.915 ;
        RECT 12.005 -22.375 12.330 -21.915 ;
        RECT 14.045 -22.375 14.315 -21.915 ;
        RECT 16.105 -22.375 16.430 -21.915 ;
        RECT -7.410 -22.545 -3.730 -22.375 ;
        RECT -3.310 -22.545 0.370 -22.375 ;
        RECT 0.790 -22.545 4.470 -22.375 ;
        RECT 5.190 -22.545 8.870 -22.375 ;
        RECT 9.290 -22.545 12.970 -22.375 ;
        RECT 13.390 -22.545 17.070 -22.375 ;
        RECT 60.600 -23.075 60.930 -22.695 ;
        RECT 61.530 -23.075 61.790 -22.235 ;
        RECT 62.150 -22.850 62.450 -22.350 ;
        RECT 60.040 -23.245 61.880 -23.075 ;
        RECT -6.850 -26.375 -6.520 -25.995 ;
        RECT -5.920 -26.375 -5.660 -25.535 ;
        RECT -5.400 -26.100 -5.000 -25.600 ;
        RECT -3.095 -26.375 -2.765 -25.995 ;
        RECT -2.155 -26.375 -1.905 -25.915 ;
        RECT -0.210 -26.375 0.160 -25.875 ;
        RECT 1.975 -26.375 2.185 -25.845 ;
        RECT 2.945 -26.375 3.115 -25.765 ;
        RECT 5.725 -26.375 6.035 -25.575 ;
        RECT 8.415 -26.375 8.645 -25.555 ;
        RECT 9.315 -26.375 9.525 -25.555 ;
        RECT -7.410 -26.545 -5.570 -26.375 ;
        RECT -3.610 -26.545 3.750 -26.375 ;
        RECT 5.640 -26.545 7.020 -26.375 ;
        RECT 8.290 -26.545 9.670 -26.375 ;
        RECT 59.650 -26.800 66.250 -26.300 ;
        RECT 59.650 -27.300 60.150 -26.800 ;
        RECT 67.920 -26.975 68.185 -26.515 ;
        RECT 68.855 -26.975 69.025 -26.515 ;
        RECT 69.695 -26.975 69.945 -26.510 ;
        RECT 72.905 -26.975 73.235 -26.595 ;
        RECT 73.845 -26.975 74.095 -26.515 ;
        RECT 75.790 -26.975 76.160 -26.475 ;
        RECT 77.975 -26.975 78.185 -26.445 ;
        RECT 78.945 -26.975 79.115 -26.365 ;
        RECT 67.790 -27.145 70.090 -26.975 ;
        RECT 72.390 -27.145 79.750 -26.975 ;
        RECT 64.850 -31.200 65.250 -30.700 ;
        RECT 66.115 -31.175 66.355 -30.695 ;
        RECT 66.945 -31.175 67.275 -30.695 ;
        RECT 67.785 -31.175 68.115 -30.375 ;
        RECT 68.350 -31.175 71.000 -31.000 ;
        RECT 71.505 -31.175 71.835 -30.795 ;
        RECT 72.445 -31.175 72.695 -30.715 ;
        RECT 74.390 -31.175 74.760 -30.675 ;
        RECT 76.575 -31.175 76.785 -30.645 ;
        RECT 77.550 -31.175 77.720 -30.565 ;
        RECT 78.390 -31.175 78.560 -30.660 ;
        RECT 79.380 -31.175 79.710 -30.435 ;
        RECT 80.305 -31.175 80.555 -30.355 ;
        RECT 65.590 -31.345 80.650 -31.175 ;
        RECT 68.350 -31.500 71.000 -31.345 ;
        RECT 42.750 -33.700 43.150 -33.200 ;
        RECT -9.800 -34.830 -9.400 -34.330 ;
        RECT -8.650 -35.005 -8.320 -34.625 ;
        RECT -7.720 -34.830 -7.460 -34.165 ;
        RECT -7.720 -35.005 -5.750 -34.830 ;
        RECT -5.255 -35.005 -4.925 -34.625 ;
        RECT -4.315 -35.005 -3.985 -34.625 ;
        RECT -2.160 -35.005 -1.750 -34.565 ;
        RECT -1.010 -35.005 -0.690 -34.545 ;
        RECT 0.920 -35.005 1.580 -34.525 ;
        RECT 2.710 -35.005 2.995 -34.545 ;
        RECT 3.850 -35.005 5.700 -34.880 ;
        RECT 6.260 -35.005 6.590 -34.625 ;
        RECT 7.190 -35.005 7.450 -34.165 ;
        RECT -9.210 -35.175 7.540 -35.005 ;
        RECT -7.500 -35.330 -5.750 -35.175 ;
        RECT 3.850 -35.330 5.700 -35.175 ;
        RECT 31.155 -35.850 31.325 -35.290 ;
        RECT 49.800 -35.300 50.200 -34.800 ;
        RECT 31.155 -36.180 31.705 -35.850 ;
        RECT 31.155 -36.780 31.325 -36.180 ;
        RECT 31.155 -37.040 32.165 -36.780 ;
        RECT 31.155 -37.130 31.325 -37.040 ;
        RECT 31.500 -37.850 32.000 -37.450 ;
        RECT 59.650 -38.000 60.150 -37.650 ;
        RECT 59.650 -38.500 66.250 -38.000 ;
        RECT 31.155 -38.715 31.325 -38.590 ;
        RECT 31.155 -38.945 32.145 -38.715 ;
        RECT 59.650 -38.850 60.150 -38.500 ;
        RECT 67.920 -38.675 68.185 -38.215 ;
        RECT 68.855 -38.675 69.025 -38.215 ;
        RECT 69.695 -38.675 69.945 -38.210 ;
        RECT 72.905 -38.675 73.235 -38.295 ;
        RECT 73.845 -38.675 74.095 -38.215 ;
        RECT 75.790 -38.675 76.160 -38.175 ;
        RECT 77.975 -38.675 78.185 -38.145 ;
        RECT 78.945 -38.675 79.115 -38.065 ;
        RECT 67.790 -38.845 70.090 -38.675 ;
        RECT 72.390 -38.845 79.750 -38.675 ;
        RECT -9.750 -40.030 -9.350 -39.530 ;
        RECT -8.935 -40.215 -8.705 -39.395 ;
        RECT -8.035 -40.030 -7.825 -39.395 ;
        RECT 31.155 -39.615 31.325 -38.945 ;
        RECT 31.155 -39.825 32.145 -39.615 ;
        RECT -8.035 -40.215 -3.150 -40.030 ;
        RECT -9.060 -40.380 -3.150 -40.215 ;
        RECT -9.060 -40.385 -7.680 -40.380 ;
        RECT -3.500 -40.580 -3.150 -40.380 ;
        RECT -0.915 -40.580 -0.585 -40.295 ;
        RECT -3.500 -40.685 -0.585 -40.580 ;
        RECT -0.075 -40.685 0.255 -40.295 ;
        RECT 1.795 -40.685 2.085 -39.850 ;
        RECT 2.600 -40.530 3.100 -40.130 ;
        RECT 4.090 -40.685 4.420 -40.305 ;
        RECT 5.020 -40.685 5.280 -39.845 ;
        RECT 31.155 -39.970 31.325 -39.825 ;
        RECT -3.500 -40.855 2.170 -40.685 ;
        RECT 3.530 -40.855 5.370 -40.685 ;
        RECT -3.500 -40.930 -0.850 -40.855 ;
        RECT -6.950 -42.655 -5.650 -42.530 ;
        RECT -3.500 -42.655 -3.150 -40.930 ;
        RECT 38.300 -41.150 43.150 -40.750 ;
        RECT 40.180 -41.990 54.200 -41.820 ;
        RECT 3.900 -42.655 6.050 -42.630 ;
        RECT -8.200 -42.825 7.700 -42.655 ;
        RECT -8.055 -43.645 -7.845 -42.825 ;
        RECT -7.175 -42.980 -5.650 -42.825 ;
        RECT -7.175 -43.645 -6.945 -42.980 ;
        RECT -4.835 -43.285 -4.550 -42.825 ;
        RECT -3.420 -43.305 -2.760 -42.825 ;
        RECT -1.150 -43.285 -0.830 -42.825 ;
        RECT -0.090 -43.265 0.320 -42.825 ;
        RECT 2.145 -43.205 2.475 -42.825 ;
        RECT 3.085 -43.205 3.415 -42.825 ;
        RECT 3.900 -42.980 6.210 -42.825 ;
        RECT 5.000 -43.380 5.500 -42.980 ;
        RECT 5.950 -43.665 6.210 -42.980 ;
        RECT 6.810 -43.205 7.140 -42.825 ;
        RECT 40.180 -43.150 40.350 -41.990 ;
        RECT 53.450 -42.470 53.750 -42.450 ;
        RECT 51.390 -42.820 53.750 -42.470 ;
        RECT 40.100 -43.300 40.500 -43.150 ;
        RECT 53.450 -43.300 53.750 -42.820 ;
        RECT 54.030 -43.300 54.200 -41.990 ;
        RECT 64.850 -42.900 65.250 -42.400 ;
        RECT 66.115 -42.875 66.355 -42.395 ;
        RECT 66.945 -42.875 67.275 -42.395 ;
        RECT 67.785 -42.875 68.115 -42.075 ;
        RECT 68.350 -42.875 71.000 -42.700 ;
        RECT 71.505 -42.875 71.835 -42.495 ;
        RECT 72.445 -42.875 72.695 -42.415 ;
        RECT 74.390 -42.875 74.760 -42.375 ;
        RECT 76.575 -42.875 76.785 -42.345 ;
        RECT 77.550 -42.875 77.720 -42.265 ;
        RECT 78.390 -42.875 78.560 -42.360 ;
        RECT 79.380 -42.875 79.710 -42.135 ;
        RECT 80.305 -42.875 80.555 -42.055 ;
        RECT 65.590 -43.045 80.650 -42.875 ;
        RECT 68.350 -43.200 71.000 -43.045 ;
        RECT 40.100 -43.470 54.200 -43.300 ;
        RECT 40.100 -43.550 40.500 -43.470 ;
      LAYER met1 ;
        RECT -6.900 26.700 -6.500 29.450 ;
        RECT 2.600 26.700 3.000 29.450 ;
        RECT 8.050 26.700 8.450 29.450 ;
        RECT 13.500 26.700 13.900 29.450 ;
        RECT 23.100 26.700 23.500 29.450 ;
        RECT 32.600 26.700 33.000 29.450 ;
        RECT 38.050 26.700 38.450 29.450 ;
        RECT 43.500 26.700 43.900 29.450 ;
        RECT 53.100 26.700 53.500 29.450 ;
        RECT 62.600 26.700 63.000 29.450 ;
        RECT 68.050 26.700 68.450 29.450 ;
        RECT 73.500 26.700 73.900 29.450 ;
        RECT -6.900 26.200 73.900 26.700 ;
        RECT 18.100 19.100 18.500 19.250 ;
        RECT 21.050 19.100 21.550 26.200 ;
        RECT 31.900 23.150 32.400 26.200 ;
        RECT 31.050 23.080 32.400 23.150 ;
        RECT 29.125 22.700 32.400 23.080 ;
        RECT 31.050 22.600 32.400 22.700 ;
        RECT 18.100 18.800 21.550 19.100 ;
        RECT 18.100 18.750 18.500 18.800 ;
        RECT 15.540 18.450 17.840 18.630 ;
        RECT 21.050 18.450 21.550 18.800 ;
        RECT 15.540 18.150 21.550 18.450 ;
        RECT 31.900 20.850 32.400 22.600 ;
        RECT 73.400 20.850 73.900 26.200 ;
        RECT 31.900 20.350 82.700 20.850 ;
        RECT 31.900 17.600 32.300 20.350 ;
        RECT 37.350 17.600 37.750 20.350 ;
        RECT 42.800 17.600 43.200 20.350 ;
        RECT 52.300 17.600 52.700 20.350 ;
        RECT 61.900 17.600 62.300 20.350 ;
        RECT 67.350 17.600 67.750 20.350 ;
        RECT 72.800 17.600 73.200 20.350 ;
        RECT 82.300 17.600 82.700 20.350 ;
        RECT -9.800 -3.180 -9.400 -2.680 ;
        RECT -9.800 -3.200 -9.100 -3.180 ;
        RECT -9.800 -3.680 -7.370 -3.200 ;
        RECT -5.770 -3.680 3.890 -3.200 ;
        RECT 5.700 -3.680 7.540 -3.200 ;
        RECT 34.600 -3.500 35.000 -3.000 ;
        RECT 39.300 -3.500 39.700 -3.000 ;
        RECT 42.400 -3.500 42.800 -3.000 ;
        RECT 45.500 -3.500 45.900 -3.000 ;
        RECT 50.200 -3.500 50.600 -3.000 ;
        RECT 54.900 -3.500 55.300 -3.000 ;
        RECT 58.000 -3.500 58.400 -3.000 ;
        RECT 61.100 -3.500 61.500 -3.000 ;
        RECT 65.800 -3.500 66.200 -3.000 ;
        RECT 70.500 -3.500 70.900 -3.000 ;
        RECT 73.600 -3.500 74.000 -3.000 ;
        RECT 76.700 -3.500 77.100 -3.000 ;
        RECT -9.750 -8.380 -9.350 -7.880 ;
        RECT -9.750 -8.410 -9.050 -8.380 ;
        RECT -9.750 -8.890 -7.680 -8.410 ;
        RECT -3.500 -8.730 -3.150 -3.680 ;
        RECT 49.050 -8.350 49.450 -7.800 ;
        RECT 2.600 -8.880 3.100 -8.480 ;
        RECT 47.600 -8.750 50.000 -8.350 ;
        RECT 91.950 -8.750 93.050 -8.250 ;
        RECT -9.750 -8.930 -9.050 -8.890 ;
        RECT -1.050 -9.360 5.370 -8.880 ;
        RECT 2.150 -9.380 3.550 -9.360 ;
        RECT 41.890 -9.550 42.200 -9.070 ;
        RECT 42.440 -9.550 44.740 -9.520 ;
        RECT 47.600 -9.550 48.100 -8.750 ;
        RECT 41.850 -10.000 48.100 -9.550 ;
        RECT 52.950 -10.100 53.350 -9.600 ;
        RECT 56.050 -10.100 56.450 -9.600 ;
        RECT 59.150 -10.100 59.550 -9.600 ;
        RECT 63.850 -10.100 64.250 -9.600 ;
        RECT 68.550 -10.100 68.950 -9.600 ;
        RECT 71.650 -10.100 72.050 -9.600 ;
        RECT 74.750 -10.100 75.150 -9.600 ;
        RECT 79.450 -10.100 79.850 -9.600 ;
        RECT -8.200 -11.330 -6.820 -10.850 ;
        RECT -5.730 -11.330 3.930 -10.850 ;
        RECT 5.860 -11.330 7.700 -10.850 ;
        RECT 12.000 -11.150 13.700 -10.650 ;
        RECT 5.000 -11.730 5.500 -11.330 ;
        RECT 11.800 -17.400 13.800 -11.150 ;
        RECT 4.650 -22.200 4.960 -21.710 ;
        RECT -3.750 -22.220 -3.300 -22.200 ;
        RECT 0.350 -22.220 0.800 -22.200 ;
        RECT 4.450 -22.220 5.200 -22.200 ;
        RECT 8.850 -22.220 9.300 -22.200 ;
        RECT 12.950 -22.220 13.400 -22.200 ;
        RECT -7.410 -22.700 17.070 -22.220 ;
        RECT -5.400 -26.200 -5.000 -25.600 ;
        RECT 12.410 -26.200 12.885 -22.700 ;
        RECT 60.040 -22.950 61.880 -22.920 ;
        RECT 62.150 -22.950 62.450 -22.350 ;
        RECT -5.600 -26.220 -3.600 -26.200 ;
        RECT 3.750 -26.220 5.650 -26.200 ;
        RECT 7.000 -26.220 8.300 -26.200 ;
        RECT 9.600 -26.220 12.885 -26.200 ;
        RECT -7.410 -26.700 12.885 -26.220 ;
        RECT 59.650 -23.400 62.450 -22.950 ;
        RECT 59.650 -26.300 60.150 -23.400 ;
        RECT -7.400 -27.900 -5.400 -26.700 ;
        RECT -0.450 -27.900 1.550 -26.700 ;
        RECT 59.650 -26.800 60.650 -26.300 ;
        RECT 65.850 -26.800 66.250 -26.300 ;
        RECT 59.650 -30.700 60.150 -26.800 ;
        RECT 67.790 -26.950 70.090 -26.820 ;
        RECT 72.390 -26.900 79.750 -26.820 ;
        RECT 72.390 -26.950 84.500 -26.900 ;
        RECT 67.790 -27.300 84.500 -26.950 ;
        RECT 59.650 -31.050 65.250 -30.700 ;
        RECT 65.590 -31.050 68.350 -31.020 ;
        RECT 59.650 -31.200 68.350 -31.050 ;
        RECT -9.800 -34.830 -9.400 -34.330 ;
        RECT -9.800 -34.850 -9.100 -34.830 ;
        RECT -9.800 -35.330 -7.370 -34.850 ;
        RECT -5.770 -35.330 3.890 -34.850 ;
        RECT 5.700 -35.330 7.540 -34.850 ;
        RECT -9.800 -35.850 -7.400 -35.330 ;
        RECT -9.750 -40.030 -9.350 -39.530 ;
        RECT -9.750 -40.060 -9.050 -40.030 ;
        RECT -9.750 -40.540 -7.680 -40.060 ;
        RECT -3.500 -40.380 -3.150 -35.330 ;
        RECT 31.000 -37.100 31.480 -35.290 ;
        RECT 31.000 -37.450 31.500 -37.100 ;
        RECT 42.750 -37.200 43.150 -33.200 ;
        RECT 49.800 -37.200 50.200 -34.800 ;
        RECT 31.000 -37.850 32.000 -37.450 ;
        RECT 42.750 -37.600 50.200 -37.200 ;
        RECT 31.000 -38.600 31.500 -37.850 ;
        RECT 31.000 -39.970 31.480 -38.600 ;
        RECT 2.600 -40.530 3.100 -40.130 ;
        RECT -9.750 -40.580 -9.050 -40.540 ;
        RECT -1.050 -41.010 5.370 -40.530 ;
        RECT 2.150 -41.030 3.550 -41.010 ;
        RECT -8.200 -42.980 -6.820 -42.500 ;
        RECT -5.730 -42.980 3.930 -42.500 ;
        RECT 5.860 -42.980 7.700 -42.500 ;
        RECT 5.000 -43.380 5.500 -42.980 ;
        RECT 31.050 -43.150 31.450 -39.970 ;
        RECT 38.300 -43.150 38.700 -40.750 ;
        RECT 42.750 -41.150 43.150 -37.600 ;
        RECT 59.650 -42.400 60.150 -31.200 ;
        RECT 64.850 -31.500 68.350 -31.200 ;
        RECT 70.990 -31.050 80.650 -31.020 ;
        RECT 84.050 -31.050 84.500 -27.300 ;
        RECT 70.990 -31.500 84.500 -31.050 ;
        RECT 65.850 -38.500 66.250 -38.000 ;
        RECT 67.790 -38.650 70.090 -38.520 ;
        RECT 72.390 -38.600 79.750 -38.520 ;
        RECT 72.390 -38.650 84.500 -38.600 ;
        RECT 67.790 -39.000 84.500 -38.650 ;
        RECT 51.415 -42.770 53.520 -42.520 ;
        RECT 59.650 -42.750 65.250 -42.400 ;
        RECT 65.590 -42.750 68.350 -42.720 ;
        RECT 59.650 -42.900 68.350 -42.750 ;
        RECT 31.050 -43.550 40.500 -43.150 ;
        RECT 40.000 -47.800 40.500 -43.550 ;
        RECT 59.650 -47.800 60.150 -42.900 ;
        RECT 64.850 -43.200 68.350 -42.900 ;
        RECT 70.990 -42.750 80.650 -42.720 ;
        RECT 84.050 -42.750 84.500 -39.000 ;
        RECT 70.990 -43.200 84.500 -42.750 ;
        RECT 92.550 -47.800 93.050 -8.750 ;
        RECT 40.000 -48.300 93.050 -47.800 ;
      LAYER met2 ;
        RECT 73.400 21.150 74.950 23.150 ;
        RECT 92.550 -11.750 93.950 -9.750 ;
        RECT 11.800 -17.400 13.800 -15.400 ;
        RECT -7.400 -29.350 -5.400 -27.350 ;
        RECT -0.450 -29.350 1.550 -27.350 ;
        RECT -9.800 -36.600 -7.400 -35.300 ;
        RECT 92.550 -36.700 93.800 -34.700 ;
        RECT 40.000 -49.000 41.950 -47.800 ;
        RECT 80.350 -49.000 82.300 -47.800 ;
      LAYER met3 ;
        RECT -20.740 49.380 106.100 52.100 ;
        RECT 73.400 21.150 106.050 23.150 ;
        RECT 92.550 -11.750 106.050 -9.750 ;
        RECT -20.650 -17.400 13.800 -15.400 ;
        RECT -20.650 -29.350 1.550 -27.350 ;
        RECT -20.650 -36.600 -7.400 -35.150 ;
        RECT -20.650 -37.150 -18.650 -36.600 ;
        RECT 92.550 -36.700 106.050 -34.700 ;
        RECT 40.000 -49.550 41.950 -48.300 ;
        RECT 80.350 -49.700 82.300 -48.300 ;
        RECT -20.740 -59.500 106.100 -56.780 ;
      LAYER met4 ;
        RECT -20.740 -59.500 -18.020 52.100 ;
        RECT 103.380 49.300 106.100 52.100 ;
        RECT 103.400 23.200 106.100 49.300 ;
        RECT 103.380 21.100 106.100 23.200 ;
        RECT 103.400 -9.700 106.100 21.100 ;
        RECT 103.380 -11.800 106.100 -9.700 ;
        RECT 103.400 -34.700 106.100 -11.800 ;
        RECT 103.380 -36.700 106.100 -34.700 ;
        RECT 40.000 -59.350 41.950 -47.750 ;
        RECT 80.350 -59.350 82.300 -47.800 ;
        RECT 103.400 -56.700 106.100 -36.700 ;
        RECT 103.380 -59.500 106.100 -56.700 ;
    END
  END GND
  OBS
      LAYER nwell ;
        RECT 34.400 -0.750 81.200 3.050 ;
        RECT 48.850 -16.150 80.050 -12.350 ;
        RECT 46.650 -28.250 50.850 -25.650 ;
        RECT 52.150 -28.300 54.550 -25.700 ;
      LAYER pwell ;
        RECT 80.650 -31.200 82.300 -30.250 ;
      LAYER nwell ;
        RECT 37.750 -37.500 41.050 -32.700 ;
        RECT 51.600 -37.550 54.900 -32.750 ;
      LAYER pwell ;
        RECT 80.650 -42.900 82.300 -41.950 ;
      LAYER li1 ;
        RECT -5.000 33.200 -3.800 33.850 ;
        RECT -6.200 28.100 -5.800 33.000 ;
        RECT -2.150 32.650 -1.750 39.050 ;
        RECT -1.300 33.200 -0.100 33.850 ;
        RECT 4.850 33.750 6.050 33.850 ;
        RECT 0.700 33.250 6.050 33.750 ;
        RECT 0.700 32.650 1.200 33.250 ;
        RECT 4.850 33.200 6.050 33.250 ;
        RECT 7.350 33.800 7.750 39.050 ;
        RECT 9.700 33.800 10.900 33.850 ;
        RECT 7.350 33.300 10.900 33.800 ;
        RECT -2.150 32.150 1.200 32.650 ;
        RECT -2.150 29.000 -1.750 32.150 ;
        RECT 1.900 28.100 2.300 33.000 ;
        RECT 3.300 28.100 3.700 33.000 ;
        RECT 7.350 29.000 7.750 33.300 ;
        RECT 9.700 33.200 10.900 33.300 ;
        RECT 8.750 28.100 9.150 33.000 ;
        RECT 12.800 29.000 13.200 39.050 ;
        RECT 15.400 33.200 16.600 33.850 ;
        RECT 14.200 28.100 14.600 33.000 ;
        RECT 18.250 29.000 18.650 39.050 ;
        RECT 19.100 33.200 20.300 33.850 ;
        RECT 25.000 33.200 26.200 33.850 ;
        RECT 22.300 28.100 22.700 33.000 ;
        RECT 23.800 28.100 24.200 33.000 ;
        RECT 27.850 32.650 28.250 39.050 ;
        RECT 28.700 33.200 29.900 33.850 ;
        RECT 34.850 33.750 36.050 33.850 ;
        RECT 30.700 33.250 36.050 33.750 ;
        RECT 30.700 32.650 31.200 33.250 ;
        RECT 34.850 33.200 36.050 33.250 ;
        RECT 37.350 33.800 37.750 39.050 ;
        RECT 39.700 33.800 40.900 33.850 ;
        RECT 37.350 33.300 40.900 33.800 ;
        RECT 27.850 32.150 31.200 32.650 ;
        RECT 27.850 29.000 28.250 32.150 ;
        RECT 31.900 28.100 32.300 33.000 ;
        RECT 33.300 28.100 33.700 33.000 ;
        RECT 37.350 29.000 37.750 33.300 ;
        RECT 39.700 33.200 40.900 33.300 ;
        RECT 38.750 28.100 39.150 33.000 ;
        RECT 42.800 29.000 43.200 39.050 ;
        RECT 45.400 33.200 46.600 33.850 ;
        RECT 44.200 28.100 44.600 33.000 ;
        RECT 48.250 29.000 48.650 39.050 ;
        RECT 49.100 33.200 50.300 33.850 ;
        RECT 55.000 33.200 56.200 33.850 ;
        RECT 52.300 28.100 52.700 33.000 ;
        RECT 53.800 28.100 54.200 33.000 ;
        RECT 57.850 32.650 58.250 39.050 ;
        RECT 58.700 33.200 59.900 33.850 ;
        RECT 64.850 33.750 66.050 33.850 ;
        RECT 60.700 33.250 66.050 33.750 ;
        RECT 60.700 32.650 61.200 33.250 ;
        RECT 64.850 33.200 66.050 33.250 ;
        RECT 67.350 33.800 67.750 39.050 ;
        RECT 69.700 33.800 70.900 33.850 ;
        RECT 67.350 33.300 70.900 33.800 ;
        RECT 57.850 32.150 61.200 32.650 ;
        RECT 57.850 29.000 58.250 32.150 ;
        RECT 61.900 28.100 62.300 33.000 ;
        RECT 63.300 28.100 63.700 33.000 ;
        RECT 67.350 29.000 67.750 33.300 ;
        RECT 69.700 33.200 70.900 33.300 ;
        RECT 68.750 28.100 69.150 33.000 ;
        RECT 72.800 29.000 73.200 39.050 ;
        RECT 75.400 33.200 76.600 33.850 ;
        RECT 74.200 28.100 74.600 33.000 ;
        RECT 78.250 29.000 78.650 39.050 ;
        RECT 79.100 33.200 80.300 33.850 ;
        RECT 82.300 28.100 82.700 33.000 ;
        RECT -6.200 27.700 82.700 28.100 ;
        RECT 23.850 24.650 24.350 27.700 ;
        RECT 24.750 24.650 25.200 24.700 ;
        RECT 23.850 24.600 25.200 24.650 ;
        RECT 23.850 24.280 27.015 24.600 ;
        RECT 23.850 24.250 25.200 24.280 ;
        RECT 23.850 23.200 24.350 24.250 ;
        RECT 24.750 24.200 25.200 24.250 ;
        RECT 23.850 23.130 25.100 23.200 ;
        RECT 23.850 23.050 25.200 23.130 ;
        RECT 23.850 22.730 27.015 23.050 ;
        RECT 23.850 22.650 25.200 22.730 ;
        RECT 23.850 22.600 25.100 22.650 ;
        RECT 15.625 20.455 15.885 20.855 ;
        RECT 17.160 20.515 17.755 20.855 ;
        RECT 15.625 20.285 16.990 20.455 ;
        RECT 16.255 19.215 16.990 20.285 ;
        RECT 15.625 19.045 16.990 19.215 ;
        RECT 17.160 19.195 17.335 20.515 ;
        RECT 23.850 19.350 24.350 22.600 ;
        RECT 81.500 19.350 82.000 27.700 ;
        RECT 15.625 18.645 15.885 19.045 ;
        RECT 17.160 18.645 17.755 19.195 ;
        RECT 23.100 18.950 82.000 19.350 ;
        RECT 23.100 14.050 23.500 18.950 ;
        RECT 25.500 13.200 26.700 13.850 ;
        RECT 27.150 8.000 27.550 18.050 ;
        RECT 31.200 14.050 31.600 18.950 ;
        RECT 29.200 13.200 30.400 13.850 ;
        RECT 32.600 8.000 33.000 18.050 ;
        RECT 36.650 14.050 37.050 18.950 ;
        RECT 34.900 13.750 36.100 13.850 ;
        RECT 38.050 13.750 38.450 18.050 ;
        RECT 42.100 14.050 42.500 18.950 ;
        RECT 43.500 14.050 43.900 18.950 ;
        RECT 47.550 14.900 47.950 18.050 ;
        RECT 44.600 14.400 47.950 14.900 ;
        RECT 34.900 13.250 38.450 13.750 ;
        RECT 34.900 13.200 36.100 13.250 ;
        RECT 38.050 8.000 38.450 13.250 ;
        RECT 39.750 13.800 40.950 13.850 ;
        RECT 44.600 13.800 45.100 14.400 ;
        RECT 39.750 13.300 45.100 13.800 ;
        RECT 39.750 13.200 40.950 13.300 ;
        RECT 45.900 13.200 47.100 13.850 ;
        RECT 47.550 8.000 47.950 14.400 ;
        RECT 51.600 14.050 52.000 18.950 ;
        RECT 53.100 14.050 53.500 18.950 ;
        RECT 49.600 13.200 50.800 13.850 ;
        RECT 55.500 13.200 56.700 13.850 ;
        RECT 57.150 8.000 57.550 18.050 ;
        RECT 61.200 14.050 61.600 18.950 ;
        RECT 59.200 13.200 60.400 13.850 ;
        RECT 62.600 8.000 63.000 18.050 ;
        RECT 66.650 14.050 67.050 18.950 ;
        RECT 64.900 13.750 66.100 13.850 ;
        RECT 68.050 13.750 68.450 18.050 ;
        RECT 72.100 14.050 72.500 18.950 ;
        RECT 73.500 14.050 73.900 18.950 ;
        RECT 77.550 14.900 77.950 18.050 ;
        RECT 74.600 14.400 77.950 14.900 ;
        RECT 64.900 13.250 68.450 13.750 ;
        RECT 64.900 13.200 66.100 13.250 ;
        RECT 68.050 8.000 68.450 13.250 ;
        RECT 69.750 13.800 70.950 13.850 ;
        RECT 74.600 13.800 75.100 14.400 ;
        RECT 69.750 13.300 75.100 13.800 ;
        RECT 69.750 13.200 70.950 13.300 ;
        RECT 75.900 13.200 77.100 13.850 ;
        RECT 77.550 8.000 77.950 14.400 ;
        RECT 81.600 14.050 82.000 18.950 ;
        RECT 79.600 13.200 80.800 13.850 ;
        RECT 34.600 3.550 81.000 3.950 ;
        RECT 34.600 2.200 35.000 3.550 ;
        RECT 35.300 -0.350 35.700 3.550 ;
        RECT -9.035 -1.735 -8.865 -0.975 ;
        RECT -9.035 -1.905 -8.320 -1.735 ;
        RECT -8.150 -1.880 -7.895 -0.975 ;
        RECT -5.595 -1.475 -5.425 -0.975 ;
        RECT -5.595 -1.645 -4.930 -1.475 ;
        RECT -10.100 -2.430 -8.750 -2.080 ;
        RECT -8.490 -2.115 -8.320 -1.905 ;
        RECT -9.125 -2.455 -8.770 -2.430 ;
        RECT -8.490 -2.445 -8.235 -2.115 ;
        RECT -8.065 -2.130 -7.895 -1.880 ;
        RECT -5.680 -2.130 -5.330 -1.815 ;
        RECT -8.065 -2.330 -5.330 -2.130 ;
        RECT -8.490 -2.635 -8.320 -2.445 ;
        RECT -8.065 -2.610 -7.895 -2.330 ;
        RECT -5.680 -2.465 -5.330 -2.330 ;
        RECT -9.035 -2.805 -8.320 -2.635 ;
        RECT -9.035 -3.185 -8.865 -2.805 ;
        RECT -8.150 -3.185 -7.895 -2.610 ;
        RECT -5.160 -2.635 -4.930 -1.645 ;
        RECT -5.595 -2.805 -4.930 -2.635 ;
        RECT -5.595 -3.095 -5.425 -2.805 ;
        RECT -4.755 -3.095 -4.530 -0.975 ;
        RECT -3.815 -1.475 -3.645 -0.975 ;
        RECT -3.410 -1.190 -2.580 -1.020 ;
        RECT -4.340 -1.645 -3.645 -1.475 ;
        RECT -4.340 -2.615 -4.170 -1.645 ;
        RECT -4.000 -2.435 -3.590 -1.815 ;
        RECT -3.420 -1.865 -2.920 -1.485 ;
        RECT -4.340 -2.805 -3.645 -2.615 ;
        RECT -3.420 -2.735 -3.200 -1.865 ;
        RECT -2.750 -2.035 -2.580 -1.190 ;
        RECT -1.780 -1.355 -1.610 -1.065 ;
        RECT -0.640 -1.275 -0.010 -1.025 ;
        RECT -0.180 -1.355 -0.010 -1.275 ;
        RECT 0.790 -1.355 1.030 -1.065 ;
        RECT -2.410 -1.605 -1.040 -1.355 ;
        RECT -2.410 -1.865 -2.160 -1.605 ;
        RECT -1.650 -2.035 -1.400 -1.875 ;
        RECT -2.750 -2.205 -1.400 -2.035 ;
        RECT -2.750 -2.245 -2.330 -2.205 ;
        RECT -3.020 -2.795 -2.670 -2.425 ;
        RECT -3.815 -3.135 -3.645 -2.805 ;
        RECT -2.500 -2.975 -2.330 -2.245 ;
        RECT -1.230 -2.375 -1.040 -1.605 ;
        RECT -2.160 -2.705 -1.750 -2.375 ;
        RECT -3.345 -3.175 -2.330 -2.975 ;
        RECT -1.460 -2.715 -1.040 -2.375 ;
        RECT -0.870 -1.785 -0.350 -1.475 ;
        RECT -0.180 -1.525 1.030 -1.355 ;
        RECT -0.870 -2.545 -0.700 -1.785 ;
        RECT -0.530 -2.375 -0.350 -1.965 ;
        RECT -0.180 -2.035 -0.010 -1.525 ;
        RECT 1.760 -1.675 1.930 -1.065 ;
        RECT 2.200 -1.525 2.530 -1.015 ;
        RECT 1.760 -1.695 2.080 -1.675 ;
        RECT 0.160 -1.865 2.080 -1.695 ;
        RECT -0.180 -2.205 1.720 -2.035 ;
        RECT 0.050 -2.545 0.380 -2.425 ;
        RECT -0.870 -2.715 0.380 -2.545 ;
        RECT -1.460 -3.145 -1.210 -2.715 ;
        RECT 0.550 -2.965 0.720 -2.205 ;
        RECT 1.390 -2.265 1.720 -2.205 ;
        RECT 0.910 -2.435 1.240 -2.375 ;
        RECT 0.910 -2.705 1.570 -2.435 ;
        RECT 1.890 -2.760 2.080 -1.865 ;
        RECT -0.130 -3.135 0.720 -2.965 ;
        RECT 1.760 -3.090 2.080 -2.760 ;
        RECT 2.280 -2.115 2.530 -1.525 ;
        RECT 3.175 -1.785 3.430 -1.115 ;
        RECT 3.250 -2.080 3.430 -1.785 ;
        RECT 5.875 -1.735 6.045 -0.975 ;
        RECT 5.875 -1.905 6.590 -1.735 ;
        RECT 6.760 -1.880 7.015 -0.975 ;
        RECT 35.950 -1.150 36.400 -0.700 ;
        RECT 3.250 -2.085 5.800 -2.080 ;
        RECT 2.280 -2.445 3.080 -2.115 ;
        RECT 2.280 -3.095 2.530 -2.445 ;
        RECT 3.250 -2.455 6.140 -2.085 ;
        RECT 6.420 -2.115 6.590 -1.905 ;
        RECT 6.420 -2.445 6.675 -2.115 ;
        RECT 3.250 -2.480 5.800 -2.455 ;
        RECT 3.250 -2.645 3.430 -2.480 ;
        RECT 6.420 -2.635 6.590 -2.445 ;
        RECT 6.845 -2.610 7.015 -1.880 ;
        RECT 3.175 -3.175 3.430 -2.645 ;
        RECT 5.875 -2.805 6.590 -2.635 ;
        RECT 5.875 -3.185 6.045 -2.805 ;
        RECT 6.760 -3.185 7.015 -2.610 ;
        RECT 36.900 -3.450 37.300 2.650 ;
        RECT 38.500 -0.350 38.900 3.550 ;
        RECT 39.300 2.600 39.700 3.550 ;
        RECT 40.000 2.600 40.400 2.650 ;
        RECT 39.300 2.100 40.400 2.600 ;
        RECT 40.000 -0.350 40.400 2.100 ;
        RECT 41.600 -0.650 42.000 2.650 ;
        RECT 42.400 2.600 42.800 3.550 ;
        RECT 43.100 2.600 43.500 2.650 ;
        RECT 42.400 2.100 43.500 2.600 ;
        RECT 43.100 -0.350 43.500 2.100 ;
        RECT 37.550 -1.150 38.000 -0.700 ;
        RECT 40.400 -1.150 41.350 -0.650 ;
        RECT 41.600 -1.150 44.450 -0.650 ;
        RECT 41.600 -3.450 42.000 -1.150 ;
        RECT 44.700 -3.450 45.100 2.650 ;
        RECT 45.500 2.200 45.900 3.550 ;
        RECT 46.200 -0.350 46.600 3.550 ;
        RECT 46.850 -1.150 47.300 -0.700 ;
        RECT 47.800 -3.450 48.200 2.650 ;
        RECT 49.400 -0.350 49.800 3.550 ;
        RECT 50.200 2.200 50.600 3.550 ;
        RECT 50.900 -0.350 51.300 3.550 ;
        RECT 48.450 -1.150 48.900 -0.700 ;
        RECT 51.550 -1.150 52.000 -0.700 ;
        RECT 52.500 -3.450 52.900 2.650 ;
        RECT 54.100 -0.350 54.500 3.550 ;
        RECT 54.900 2.600 55.300 3.550 ;
        RECT 55.600 2.600 56.000 2.650 ;
        RECT 54.900 2.100 56.000 2.600 ;
        RECT 55.600 -0.350 56.000 2.100 ;
        RECT 57.200 -0.650 57.600 2.650 ;
        RECT 58.000 2.600 58.400 3.550 ;
        RECT 58.700 2.600 59.100 2.650 ;
        RECT 58.000 2.100 59.100 2.600 ;
        RECT 58.700 -0.350 59.100 2.100 ;
        RECT 53.150 -1.150 53.600 -0.700 ;
        RECT 56.000 -1.150 56.950 -0.650 ;
        RECT 57.200 -1.150 60.050 -0.650 ;
        RECT 57.200 -3.450 57.600 -1.150 ;
        RECT 60.300 -3.450 60.700 2.650 ;
        RECT 61.100 2.200 61.500 3.550 ;
        RECT 61.800 -0.350 62.200 3.550 ;
        RECT 62.450 -1.150 62.900 -0.700 ;
        RECT 63.400 -3.450 63.800 2.650 ;
        RECT 65.000 -0.350 65.400 3.550 ;
        RECT 65.800 2.200 66.200 3.550 ;
        RECT 66.500 -0.350 66.900 3.550 ;
        RECT 64.050 -1.150 64.500 -0.700 ;
        RECT 67.150 -1.150 67.600 -0.700 ;
        RECT 68.100 -3.450 68.500 2.650 ;
        RECT 69.700 -0.350 70.100 3.550 ;
        RECT 70.500 2.600 70.900 3.550 ;
        RECT 71.200 2.600 71.600 2.650 ;
        RECT 70.500 2.100 71.600 2.600 ;
        RECT 71.200 -0.350 71.600 2.100 ;
        RECT 72.800 -0.650 73.200 2.650 ;
        RECT 73.600 2.600 74.000 3.550 ;
        RECT 74.300 2.600 74.700 2.650 ;
        RECT 73.600 2.100 74.700 2.600 ;
        RECT 74.300 -0.350 74.700 2.100 ;
        RECT 68.750 -1.150 69.200 -0.700 ;
        RECT 71.600 -1.150 72.550 -0.650 ;
        RECT 72.800 -1.150 75.650 -0.650 ;
        RECT 72.800 -3.450 73.200 -1.150 ;
        RECT 75.900 -3.450 76.300 2.650 ;
        RECT 76.700 2.200 77.100 3.550 ;
        RECT 77.400 -0.350 77.800 3.550 ;
        RECT 78.050 -1.150 78.500 -0.700 ;
        RECT 79.000 -3.450 79.400 2.650 ;
        RECT 80.600 -0.350 81.000 3.550 ;
        RECT 79.650 -1.150 80.100 -0.700 ;
        RECT -8.535 -7.165 -8.205 -6.185 ;
        RECT -8.455 -7.380 -8.205 -7.165 ;
        RECT -0.965 -7.335 -0.585 -6.655 ;
        RECT 0.345 -7.165 0.675 -6.655 ;
        RECT 1.185 -7.165 1.585 -6.655 ;
        RECT 0.345 -7.335 1.585 -7.165 ;
        RECT -8.455 -7.550 -8.200 -7.380 ;
        RECT -8.455 -7.765 -8.205 -7.550 ;
        RECT -8.535 -8.395 -8.205 -7.765 ;
        RECT -0.965 -8.295 -0.795 -7.335 ;
        RECT -0.625 -7.675 0.680 -7.505 ;
        RECT 1.765 -7.585 2.085 -6.655 ;
        RECT 3.705 -7.415 3.875 -6.655 ;
        RECT 3.705 -7.585 4.420 -7.415 ;
        RECT 4.590 -7.560 4.845 -6.655 ;
        RECT -0.625 -8.125 -0.380 -7.675 ;
        RECT -0.210 -8.045 0.340 -7.845 ;
        RECT 0.510 -7.875 0.680 -7.675 ;
        RECT 1.455 -7.730 2.085 -7.585 ;
        RECT 1.455 -7.780 3.300 -7.730 ;
        RECT 3.615 -7.780 3.970 -7.765 ;
        RECT 0.510 -8.045 0.885 -7.875 ;
        RECT 1.055 -8.295 1.285 -7.795 ;
        RECT -0.965 -8.465 1.285 -8.295 ;
        RECT 1.455 -7.980 3.970 -7.780 ;
        RECT -0.415 -8.785 -0.245 -8.465 ;
        RECT 1.455 -8.635 1.625 -7.980 ;
        RECT 3.615 -8.135 3.970 -7.980 ;
        RECT 4.250 -7.795 4.420 -7.585 ;
        RECT 4.250 -8.125 4.505 -7.795 ;
        RECT 4.250 -8.315 4.420 -8.125 ;
        RECT 4.675 -8.290 4.845 -7.560 ;
        RECT 42.525 -7.695 42.785 -7.295 ;
        RECT 44.060 -7.300 44.655 -7.295 ;
        RECT 44.060 -7.600 46.950 -7.300 ;
        RECT 44.060 -7.635 44.655 -7.600 ;
        RECT 5.650 -8.100 30.550 -7.700 ;
        RECT 42.525 -7.865 43.890 -7.695 ;
        RECT 0.670 -8.805 1.625 -8.635 ;
        RECT 3.705 -8.485 4.420 -8.315 ;
        RECT 3.705 -8.865 3.875 -8.485 ;
        RECT 4.590 -8.865 4.845 -8.290 ;
        RECT 30.150 -8.500 30.550 -8.100 ;
        RECT 43.155 -8.935 43.890 -7.865 ;
        RECT 42.525 -9.105 43.890 -8.935 ;
        RECT 44.060 -8.955 44.235 -7.635 ;
        RECT 42.525 -9.505 42.785 -9.105 ;
        RECT 44.060 -9.505 44.655 -8.955 ;
        RECT 46.650 -10.450 46.950 -7.600 ;
        RECT 46.600 -10.850 47.000 -10.450 ;
        RECT -7.675 -11.975 -7.345 -11.345 ;
        RECT -5.270 -11.885 -5.015 -11.355 ;
        RECT -7.675 -12.575 -7.425 -11.975 ;
        RECT -7.255 -12.170 -6.925 -12.165 ;
        RECT -5.270 -12.170 -5.090 -11.885 ;
        RECT -4.370 -12.085 -4.120 -11.435 ;
        RECT -7.255 -12.410 -5.090 -12.170 ;
        RECT -7.255 -12.415 -6.925 -12.410 ;
        RECT -7.675 -13.555 -7.345 -12.575 ;
        RECT -5.270 -12.745 -5.090 -12.410 ;
        RECT -4.920 -12.415 -4.120 -12.085 ;
        RECT -5.270 -13.415 -5.015 -12.745 ;
        RECT -4.370 -13.005 -4.120 -12.415 ;
        RECT -3.920 -11.770 -3.600 -11.440 ;
        RECT -2.560 -11.565 -1.710 -11.395 ;
        RECT -3.920 -12.665 -3.730 -11.770 ;
        RECT -3.410 -12.095 -2.750 -11.825 ;
        RECT -3.080 -12.155 -2.750 -12.095 ;
        RECT -3.560 -12.325 -3.230 -12.265 ;
        RECT -2.560 -12.325 -2.390 -11.565 ;
        RECT -0.630 -11.815 -0.380 -11.385 ;
        RECT -2.220 -11.985 -0.970 -11.815 ;
        RECT -2.220 -12.105 -1.890 -11.985 ;
        RECT -3.560 -12.495 -1.660 -12.325 ;
        RECT -3.920 -12.835 -2.000 -12.665 ;
        RECT -3.920 -12.855 -3.600 -12.835 ;
        RECT -4.370 -13.515 -4.040 -13.005 ;
        RECT -3.770 -13.465 -3.600 -12.855 ;
        RECT -1.830 -13.005 -1.660 -12.495 ;
        RECT -1.490 -12.565 -1.310 -12.155 ;
        RECT -1.140 -12.745 -0.970 -11.985 ;
        RECT -2.870 -13.175 -1.660 -13.005 ;
        RECT -1.490 -13.055 -0.970 -12.745 ;
        RECT -0.800 -12.155 -0.380 -11.815 ;
        RECT 0.490 -11.555 1.505 -11.355 ;
        RECT -0.090 -12.155 0.320 -11.825 ;
        RECT -0.800 -12.925 -0.610 -12.155 ;
        RECT 0.490 -12.285 0.660 -11.555 ;
        RECT 1.805 -11.725 1.975 -11.395 ;
        RECT 0.830 -12.105 1.180 -11.735 ;
        RECT 0.490 -12.325 0.910 -12.285 ;
        RECT -0.440 -12.495 0.910 -12.325 ;
        RECT -0.440 -12.655 -0.190 -12.495 ;
        RECT 0.320 -12.925 0.570 -12.665 ;
        RECT -0.800 -13.175 0.570 -12.925 ;
        RECT -2.870 -13.465 -2.630 -13.175 ;
        RECT -1.830 -13.255 -1.660 -13.175 ;
        RECT -1.830 -13.505 -1.200 -13.255 ;
        RECT -0.230 -13.465 -0.060 -13.175 ;
        RECT 0.740 -13.340 0.910 -12.495 ;
        RECT 1.360 -12.665 1.580 -11.795 ;
        RECT 1.805 -11.915 2.500 -11.725 ;
        RECT 1.080 -13.045 1.580 -12.665 ;
        RECT 1.750 -12.715 2.160 -12.095 ;
        RECT 2.330 -12.885 2.500 -11.915 ;
        RECT 1.805 -13.055 2.500 -12.885 ;
        RECT 0.740 -13.510 1.570 -13.340 ;
        RECT 1.805 -13.555 1.975 -13.055 ;
        RECT 2.690 -13.555 2.915 -11.435 ;
        RECT 3.585 -11.725 3.755 -11.435 ;
        RECT 3.090 -11.895 3.755 -11.725 ;
        RECT 3.090 -12.885 3.320 -11.895 ;
        RECT 6.385 -11.920 6.640 -11.345 ;
        RECT 7.355 -11.725 7.525 -11.345 ;
        RECT 6.810 -11.895 7.525 -11.725 ;
        RECT 3.490 -12.080 3.840 -12.065 ;
        RECT 3.490 -12.430 5.400 -12.080 ;
        RECT 3.490 -12.715 3.840 -12.430 ;
        RECT 6.385 -12.650 6.555 -11.920 ;
        RECT 6.810 -12.085 6.980 -11.895 ;
        RECT 7.900 -12.070 19.750 -12.000 ;
        RECT 6.725 -12.415 6.980 -12.085 ;
        RECT 6.810 -12.625 6.980 -12.415 ;
        RECT 7.260 -12.450 19.750 -12.070 ;
        RECT 49.950 -12.400 50.400 -11.950 ;
        RECT 7.900 -12.500 19.750 -12.450 ;
        RECT 3.090 -13.055 3.755 -12.885 ;
        RECT 3.585 -13.555 3.755 -13.055 ;
        RECT 6.385 -13.555 6.640 -12.650 ;
        RECT 6.810 -12.795 7.525 -12.625 ;
        RECT 7.355 -13.555 7.525 -12.795 ;
        RECT 19.250 -13.000 19.750 -12.500 ;
        RECT 49.050 -16.650 49.450 -12.750 ;
        RECT 50.650 -15.750 51.050 -9.650 ;
        RECT 51.550 -12.400 52.000 -11.950 ;
        RECT 52.250 -16.650 52.650 -12.750 ;
        RECT 52.950 -16.650 53.350 -15.300 ;
        RECT 53.750 -15.750 54.150 -9.650 ;
        RECT 56.850 -11.950 57.250 -9.650 ;
        RECT 54.400 -12.450 57.250 -11.950 ;
        RECT 57.500 -12.450 58.450 -11.950 ;
        RECT 60.850 -12.400 61.300 -11.950 ;
        RECT 55.350 -15.200 55.750 -12.750 ;
        RECT 55.350 -15.700 56.450 -15.200 ;
        RECT 55.350 -15.750 55.750 -15.700 ;
        RECT 56.050 -16.650 56.450 -15.700 ;
        RECT 56.850 -15.750 57.250 -12.450 ;
        RECT 58.450 -15.200 58.850 -12.750 ;
        RECT 58.450 -15.700 59.550 -15.200 ;
        RECT 58.450 -15.750 58.850 -15.700 ;
        RECT 59.150 -16.650 59.550 -15.700 ;
        RECT 59.950 -16.650 60.350 -12.750 ;
        RECT 61.550 -15.750 61.950 -9.650 ;
        RECT 62.450 -12.400 62.900 -11.950 ;
        RECT 65.550 -12.400 66.000 -11.950 ;
        RECT 63.150 -16.650 63.550 -12.750 ;
        RECT 63.850 -16.650 64.250 -15.300 ;
        RECT 64.650 -16.650 65.050 -12.750 ;
        RECT 66.250 -15.750 66.650 -9.650 ;
        RECT 67.150 -12.400 67.600 -11.950 ;
        RECT 67.850 -16.650 68.250 -12.750 ;
        RECT 68.550 -16.650 68.950 -15.300 ;
        RECT 69.350 -15.750 69.750 -9.650 ;
        RECT 72.450 -11.950 72.850 -9.650 ;
        RECT 70.000 -12.450 72.850 -11.950 ;
        RECT 73.100 -12.450 74.050 -11.950 ;
        RECT 76.450 -12.400 76.900 -11.950 ;
        RECT 70.950 -15.200 71.350 -12.750 ;
        RECT 70.950 -15.700 72.050 -15.200 ;
        RECT 70.950 -15.750 71.350 -15.700 ;
        RECT 71.650 -16.650 72.050 -15.700 ;
        RECT 72.450 -15.750 72.850 -12.450 ;
        RECT 74.050 -15.200 74.450 -12.750 ;
        RECT 74.050 -15.700 75.150 -15.200 ;
        RECT 74.050 -15.750 74.450 -15.700 ;
        RECT 74.750 -16.650 75.150 -15.700 ;
        RECT 75.550 -16.650 75.950 -12.750 ;
        RECT 77.150 -15.750 77.550 -9.650 ;
        RECT 78.050 -12.400 78.500 -11.950 ;
        RECT 78.750 -16.650 79.150 -12.750 ;
        RECT 79.450 -16.650 79.850 -15.300 ;
        RECT 49.050 -17.050 79.850 -16.650 ;
        RECT -7.210 -20.455 -6.925 -19.995 ;
        RECT -7.210 -20.675 -6.255 -20.455 ;
        RECT -6.465 -21.575 -6.255 -20.675 ;
        RECT -7.210 -21.745 -6.255 -21.575 ;
        RECT -6.085 -20.845 -5.685 -19.995 ;
        RECT -5.495 -20.455 -5.215 -19.995 ;
        RECT -5.495 -20.675 -4.370 -20.455 ;
        RECT -6.085 -21.405 -4.990 -20.845 ;
        RECT -4.820 -21.135 -4.370 -20.675 ;
        RECT -4.200 -20.850 -3.815 -19.995 ;
        RECT -3.110 -20.455 -2.825 -19.995 ;
        RECT -3.110 -20.675 -2.155 -20.455 ;
        RECT -3.225 -20.850 -2.535 -20.845 ;
        RECT -4.200 -20.965 -2.535 -20.850 ;
        RECT -7.210 -22.205 -6.925 -21.745 ;
        RECT -6.085 -22.205 -5.685 -21.405 ;
        RECT -4.820 -21.465 -4.265 -21.135 ;
        RECT -4.095 -21.400 -2.535 -20.965 ;
        RECT -4.820 -21.575 -4.370 -21.465 ;
        RECT -5.495 -21.745 -4.370 -21.575 ;
        RECT -4.095 -21.635 -3.815 -21.400 ;
        RECT -3.225 -21.405 -2.535 -21.400 ;
        RECT -2.365 -21.575 -2.155 -20.675 ;
        RECT -5.495 -22.205 -5.215 -21.745 ;
        RECT -4.200 -22.205 -3.815 -21.635 ;
        RECT -3.110 -21.745 -2.155 -21.575 ;
        RECT -1.985 -20.845 -1.585 -19.995 ;
        RECT -1.395 -20.455 -1.115 -19.995 ;
        RECT -1.395 -20.675 -0.270 -20.455 ;
        RECT -1.985 -21.405 -0.890 -20.845 ;
        RECT -0.720 -21.135 -0.270 -20.675 ;
        RECT -0.100 -20.850 0.285 -19.995 ;
        RECT 0.990 -20.455 1.275 -19.995 ;
        RECT 0.990 -20.675 1.945 -20.455 ;
        RECT 0.875 -20.850 1.565 -20.845 ;
        RECT -0.100 -20.965 1.565 -20.850 ;
        RECT -3.110 -22.205 -2.825 -21.745 ;
        RECT -1.985 -22.205 -1.585 -21.405 ;
        RECT -0.720 -21.465 -0.165 -21.135 ;
        RECT 0.005 -21.400 1.565 -20.965 ;
        RECT -0.720 -21.575 -0.270 -21.465 ;
        RECT -1.395 -21.745 -0.270 -21.575 ;
        RECT 0.005 -21.635 0.285 -21.400 ;
        RECT 0.875 -21.405 1.565 -21.400 ;
        RECT 1.735 -21.575 1.945 -20.675 ;
        RECT -1.395 -22.205 -1.115 -21.745 ;
        RECT -0.100 -22.205 0.285 -21.635 ;
        RECT 0.990 -21.745 1.945 -21.575 ;
        RECT 2.115 -20.845 2.515 -19.995 ;
        RECT 2.705 -20.455 2.985 -19.995 ;
        RECT 2.705 -20.675 3.830 -20.455 ;
        RECT 2.115 -21.405 3.210 -20.845 ;
        RECT 3.380 -21.135 3.830 -20.675 ;
        RECT 4.000 -20.850 4.385 -19.995 ;
        RECT 5.390 -20.455 5.675 -19.995 ;
        RECT 5.390 -20.675 6.345 -20.455 ;
        RECT 5.275 -20.850 5.965 -20.845 ;
        RECT 4.000 -20.965 5.965 -20.850 ;
        RECT 0.990 -22.205 1.275 -21.745 ;
        RECT 2.115 -22.205 2.515 -21.405 ;
        RECT 3.380 -21.465 3.935 -21.135 ;
        RECT 4.105 -21.400 5.965 -20.965 ;
        RECT 3.380 -21.575 3.830 -21.465 ;
        RECT 2.705 -21.745 3.830 -21.575 ;
        RECT 4.105 -21.635 4.385 -21.400 ;
        RECT 5.275 -21.405 5.965 -21.400 ;
        RECT 6.135 -21.575 6.345 -20.675 ;
        RECT 2.705 -22.205 2.985 -21.745 ;
        RECT 4.000 -22.205 4.385 -21.635 ;
        RECT 5.390 -21.745 6.345 -21.575 ;
        RECT 6.515 -20.845 6.915 -19.995 ;
        RECT 7.105 -20.455 7.385 -19.995 ;
        RECT 7.105 -20.675 8.230 -20.455 ;
        RECT 6.515 -21.405 7.610 -20.845 ;
        RECT 7.780 -21.135 8.230 -20.675 ;
        RECT 8.400 -20.850 8.785 -19.995 ;
        RECT 9.490 -20.455 9.775 -19.995 ;
        RECT 9.490 -20.675 10.445 -20.455 ;
        RECT 9.375 -20.850 10.065 -20.845 ;
        RECT 8.400 -20.965 10.065 -20.850 ;
        RECT 5.390 -22.205 5.675 -21.745 ;
        RECT 6.515 -22.205 6.915 -21.405 ;
        RECT 7.780 -21.465 8.335 -21.135 ;
        RECT 8.505 -21.400 10.065 -20.965 ;
        RECT 7.780 -21.575 8.230 -21.465 ;
        RECT 7.105 -21.745 8.230 -21.575 ;
        RECT 8.505 -21.635 8.785 -21.400 ;
        RECT 9.375 -21.405 10.065 -21.400 ;
        RECT 10.235 -21.575 10.445 -20.675 ;
        RECT 7.105 -22.205 7.385 -21.745 ;
        RECT 8.400 -22.205 8.785 -21.635 ;
        RECT 9.490 -21.745 10.445 -21.575 ;
        RECT 10.615 -20.845 11.015 -19.995 ;
        RECT 11.205 -20.455 11.485 -19.995 ;
        RECT 11.205 -20.675 12.330 -20.455 ;
        RECT 10.615 -21.405 11.710 -20.845 ;
        RECT 11.880 -21.135 12.330 -20.675 ;
        RECT 12.500 -20.850 12.885 -19.995 ;
        RECT 13.590 -20.455 13.875 -19.995 ;
        RECT 13.590 -20.675 14.545 -20.455 ;
        RECT 13.475 -20.850 14.165 -20.845 ;
        RECT 12.500 -20.965 14.165 -20.850 ;
        RECT 9.490 -22.205 9.775 -21.745 ;
        RECT 10.615 -22.205 11.015 -21.405 ;
        RECT 11.880 -21.465 12.435 -21.135 ;
        RECT 12.605 -21.400 14.165 -20.965 ;
        RECT 11.880 -21.575 12.330 -21.465 ;
        RECT 11.205 -21.745 12.330 -21.575 ;
        RECT 12.605 -21.635 12.885 -21.400 ;
        RECT 13.475 -21.405 14.165 -21.400 ;
        RECT 14.335 -21.575 14.545 -20.675 ;
        RECT 11.205 -22.205 11.485 -21.745 ;
        RECT 12.500 -22.205 12.885 -21.635 ;
        RECT 13.590 -21.745 14.545 -21.575 ;
        RECT 14.715 -20.845 15.115 -19.995 ;
        RECT 15.305 -20.455 15.585 -19.995 ;
        RECT 15.305 -20.675 16.430 -20.455 ;
        RECT 14.715 -21.405 15.810 -20.845 ;
        RECT 15.980 -21.135 16.430 -20.675 ;
        RECT 16.600 -20.965 16.985 -19.995 ;
        RECT 13.590 -22.205 13.875 -21.745 ;
        RECT 14.715 -22.205 15.115 -21.405 ;
        RECT 15.980 -21.465 16.535 -21.135 ;
        RECT 15.980 -21.575 16.430 -21.465 ;
        RECT 15.305 -21.745 16.430 -21.575 ;
        RECT 16.705 -21.550 16.985 -20.965 ;
        RECT 16.705 -21.635 18.400 -21.550 ;
        RECT 15.305 -22.205 15.585 -21.745 ;
        RECT 16.600 -21.900 18.400 -21.635 ;
        RECT 16.600 -22.205 16.985 -21.900 ;
        RECT 18.050 -22.900 18.400 -21.900 ;
        RECT 7.450 -23.250 18.400 -22.900 ;
        RECT -7.235 -24.755 -7.065 -23.995 ;
        RECT -7.235 -24.925 -6.520 -24.755 ;
        RECT -6.350 -24.900 -6.095 -23.995 ;
        RECT -3.435 -24.495 -3.265 -23.995 ;
        RECT -3.435 -24.665 -2.770 -24.495 ;
        RECT -7.325 -25.475 -6.970 -25.105 ;
        RECT -6.690 -25.135 -6.520 -24.925 ;
        RECT -6.690 -25.465 -6.435 -25.135 ;
        RECT -6.690 -25.655 -6.520 -25.465 ;
        RECT -6.265 -25.630 -6.095 -24.900 ;
        RECT -7.235 -25.825 -6.520 -25.655 ;
        RECT -7.235 -26.205 -7.065 -25.825 ;
        RECT -6.350 -26.205 -6.095 -25.630 ;
        RECT -3.000 -25.655 -2.770 -24.665 ;
        RECT -3.435 -25.825 -2.770 -25.655 ;
        RECT -3.435 -26.115 -3.265 -25.825 ;
        RECT -2.595 -26.115 -2.410 -23.995 ;
        RECT -1.735 -24.420 -1.485 -23.995 ;
        RECT -1.275 -24.270 -0.170 -24.100 ;
        RECT -1.790 -24.550 -1.485 -24.420 ;
        RECT -2.240 -25.745 -1.960 -24.795 ;
        RECT -1.790 -25.655 -1.620 -24.550 ;
        RECT -1.450 -25.335 -1.210 -24.740 ;
        RECT -1.040 -24.805 -0.510 -24.440 ;
        RECT -1.040 -25.505 -0.870 -24.805 ;
        RECT -0.340 -24.885 -0.170 -24.270 ;
        RECT 0.340 -24.325 0.590 -23.995 ;
        RECT 0.815 -24.295 1.700 -24.125 ;
        RECT -0.340 -24.975 0.170 -24.885 ;
        RECT -1.790 -25.785 -1.565 -25.655 ;
        RECT -1.395 -25.725 -0.870 -25.505 ;
        RECT -0.700 -25.145 0.170 -24.975 ;
        RECT -1.735 -25.925 -1.565 -25.785 ;
        RECT -0.700 -25.925 -0.530 -25.145 ;
        RECT 0.000 -25.215 0.170 -25.145 ;
        RECT -0.320 -25.395 -0.120 -25.365 ;
        RECT 0.340 -25.395 0.510 -24.325 ;
        RECT 0.680 -25.215 0.870 -24.495 ;
        RECT -0.320 -25.695 0.510 -25.395 ;
        RECT 1.040 -25.425 1.360 -24.465 ;
        RECT -1.735 -26.095 -1.400 -25.925 ;
        RECT -1.205 -26.095 -0.530 -25.925 ;
        RECT 0.340 -25.925 0.510 -25.695 ;
        RECT 0.895 -25.755 1.360 -25.425 ;
        RECT 1.530 -25.135 1.700 -24.295 ;
        RECT 2.425 -24.555 2.765 -23.995 ;
        RECT 1.870 -24.930 2.765 -24.555 ;
        RECT 2.575 -25.135 2.765 -24.930 ;
        RECT 6.175 -24.975 6.505 -23.995 ;
        RECT 1.530 -25.465 2.405 -25.135 ;
        RECT 2.575 -25.465 3.325 -25.135 ;
        RECT 1.530 -25.925 1.700 -25.465 ;
        RECT 2.575 -25.635 2.775 -25.465 ;
        RECT 0.340 -26.095 0.745 -25.925 ;
        RECT 0.915 -26.095 1.700 -25.925 ;
        RECT 2.445 -26.160 2.775 -25.635 ;
        RECT 6.240 -25.575 6.410 -24.975 ;
        RECT 6.580 -25.150 6.915 -25.135 ;
        RECT 7.450 -25.150 7.800 -23.250 ;
        RECT 8.815 -24.975 9.145 -23.995 ;
        RECT 19.250 -24.350 19.750 -23.850 ;
        RECT 10.400 -24.850 19.750 -24.350 ;
        RECT 6.580 -25.385 7.800 -25.150 ;
        RECT 8.395 -25.385 8.725 -25.135 ;
        RECT 6.900 -25.400 7.800 -25.385 ;
        RECT 8.895 -25.575 9.145 -24.975 ;
        RECT 19.250 -25.350 19.750 -24.850 ;
        RECT 6.240 -26.205 6.935 -25.575 ;
        RECT 8.815 -26.205 9.145 -25.575 ;
        RECT 39.200 -27.850 39.600 -26.050 ;
        RECT 42.950 -27.850 43.350 -26.050 ;
        RECT 44.750 -28.600 45.150 -26.050 ;
        RECT 46.850 -28.600 47.250 -26.000 ;
        RECT 47.550 -28.600 47.950 -26.050 ;
        RECT 44.750 -29.000 47.950 -28.600 ;
        RECT 48.450 -30.550 48.850 -26.050 ;
        RECT 49.350 -27.850 49.750 -26.050 ;
        RECT 50.250 -27.850 50.650 -26.050 ;
        RECT 52.350 -26.550 52.750 -26.050 ;
        RECT 53.050 -27.900 53.450 -26.100 ;
        RECT 53.950 -27.400 54.350 -26.100 ;
        RECT 55.900 -27.400 56.400 -17.050 ;
        RECT 60.215 -21.455 60.385 -20.695 ;
        RECT 60.215 -21.625 60.930 -21.455 ;
        RECT 61.100 -21.600 61.355 -20.695 ;
        RECT 60.125 -22.175 60.480 -21.805 ;
        RECT 60.760 -21.835 60.930 -21.625 ;
        RECT 60.760 -22.165 61.015 -21.835 ;
        RECT 60.760 -22.355 60.930 -22.165 ;
        RECT 61.185 -22.330 61.355 -21.600 ;
        RECT 60.215 -22.525 60.930 -22.355 ;
        RECT 60.215 -22.905 60.385 -22.525 ;
        RECT 61.100 -22.905 61.355 -22.330 ;
        RECT 68.355 -25.395 68.685 -24.595 ;
        RECT 69.195 -25.375 69.525 -24.595 ;
        RECT 72.565 -25.095 72.735 -24.595 ;
        RECT 72.565 -25.265 73.230 -25.095 ;
        RECT 69.195 -25.395 69.960 -25.375 ;
        RECT 68.355 -25.450 69.960 -25.395 ;
        RECT 72.480 -25.450 72.830 -25.435 ;
        RECT 68.355 -25.565 72.830 -25.450 ;
        RECT 67.895 -25.985 69.525 -25.735 ;
        RECT 69.695 -25.850 72.830 -25.565 ;
        RECT 69.695 -26.155 69.960 -25.850 ;
        RECT 72.480 -26.085 72.830 -25.850 ;
        RECT 68.355 -26.335 69.960 -26.155 ;
        RECT 73.000 -26.255 73.230 -25.265 ;
        RECT 68.355 -26.805 68.685 -26.335 ;
        RECT 69.195 -26.805 69.525 -26.335 ;
        RECT 71.000 -26.750 71.550 -26.300 ;
        RECT 72.565 -26.425 73.230 -26.255 ;
        RECT 72.565 -26.715 72.735 -26.425 ;
        RECT 73.405 -26.715 73.590 -24.595 ;
        RECT 74.265 -25.020 74.515 -24.595 ;
        RECT 74.725 -24.870 75.830 -24.700 ;
        RECT 74.210 -25.150 74.515 -25.020 ;
        RECT 73.760 -26.345 74.040 -25.395 ;
        RECT 74.210 -26.255 74.380 -25.150 ;
        RECT 74.550 -25.935 74.790 -25.340 ;
        RECT 74.960 -25.405 75.490 -25.040 ;
        RECT 74.960 -26.105 75.130 -25.405 ;
        RECT 75.660 -25.485 75.830 -24.870 ;
        RECT 76.340 -24.925 76.590 -24.595 ;
        RECT 76.815 -24.895 77.700 -24.725 ;
        RECT 75.660 -25.575 76.170 -25.485 ;
        RECT 74.210 -26.385 74.435 -26.255 ;
        RECT 74.605 -26.325 75.130 -26.105 ;
        RECT 75.300 -25.745 76.170 -25.575 ;
        RECT 74.265 -26.525 74.435 -26.385 ;
        RECT 75.300 -26.525 75.470 -25.745 ;
        RECT 76.000 -25.815 76.170 -25.745 ;
        RECT 75.680 -25.995 75.880 -25.965 ;
        RECT 76.340 -25.995 76.510 -24.925 ;
        RECT 76.680 -25.815 76.870 -25.095 ;
        RECT 75.680 -26.295 76.510 -25.995 ;
        RECT 77.040 -26.025 77.360 -25.065 ;
        RECT 74.265 -26.695 74.600 -26.525 ;
        RECT 74.795 -26.695 75.470 -26.525 ;
        RECT 76.340 -26.525 76.510 -26.295 ;
        RECT 76.895 -26.355 77.360 -26.025 ;
        RECT 77.530 -25.735 77.700 -24.895 ;
        RECT 78.425 -25.155 78.765 -24.595 ;
        RECT 77.870 -25.530 78.765 -25.155 ;
        RECT 78.575 -25.735 78.765 -25.530 ;
        RECT 79.275 -25.485 79.605 -24.640 ;
        RECT 79.275 -25.565 79.665 -25.485 ;
        RECT 79.450 -25.615 79.665 -25.565 ;
        RECT 77.530 -26.065 78.405 -25.735 ;
        RECT 78.575 -26.065 79.325 -25.735 ;
        RECT 77.530 -26.525 77.700 -26.065 ;
        RECT 78.575 -26.235 78.775 -26.065 ;
        RECT 79.495 -26.195 79.665 -25.615 ;
        RECT 79.440 -26.235 79.665 -26.195 ;
        RECT 76.340 -26.695 76.745 -26.525 ;
        RECT 76.915 -26.695 77.700 -26.525 ;
        RECT 53.950 -27.900 56.400 -27.400 ;
        RECT 71.175 -27.625 71.425 -26.750 ;
        RECT 78.445 -26.760 78.775 -26.235 ;
        RECT 79.285 -26.320 79.665 -26.235 ;
        RECT 79.285 -26.755 79.615 -26.320 ;
        RECT 40.350 -31.050 52.200 -30.550 ;
        RECT 40.350 -31.550 40.850 -31.050 ;
        RECT 37.950 -32.050 40.850 -31.550 ;
        RECT -9.035 -33.385 -8.865 -32.625 ;
        RECT -9.035 -33.555 -8.320 -33.385 ;
        RECT -8.150 -33.530 -7.895 -32.625 ;
        RECT -5.595 -33.125 -5.425 -32.625 ;
        RECT -5.595 -33.295 -4.930 -33.125 ;
        RECT -11.200 -33.730 -9.150 -33.700 ;
        RECT -11.200 -34.080 -8.750 -33.730 ;
        RECT -8.490 -33.765 -8.320 -33.555 ;
        RECT -11.200 -34.100 -8.770 -34.080 ;
        RECT -11.200 -34.500 -10.800 -34.100 ;
        RECT -9.125 -34.105 -8.770 -34.100 ;
        RECT -8.490 -34.095 -8.235 -33.765 ;
        RECT -8.065 -33.780 -7.895 -33.530 ;
        RECT -5.680 -33.780 -5.330 -33.465 ;
        RECT -8.065 -33.980 -5.330 -33.780 ;
        RECT -8.490 -34.285 -8.320 -34.095 ;
        RECT -8.065 -34.260 -7.895 -33.980 ;
        RECT -5.680 -34.115 -5.330 -33.980 ;
        RECT -9.035 -34.455 -8.320 -34.285 ;
        RECT -9.035 -34.835 -8.865 -34.455 ;
        RECT -8.150 -34.835 -7.895 -34.260 ;
        RECT -5.160 -34.285 -4.930 -33.295 ;
        RECT -5.595 -34.455 -4.930 -34.285 ;
        RECT -5.595 -34.745 -5.425 -34.455 ;
        RECT -4.755 -34.745 -4.530 -32.625 ;
        RECT -3.815 -33.125 -3.645 -32.625 ;
        RECT -3.410 -32.840 -2.580 -32.670 ;
        RECT -4.340 -33.295 -3.645 -33.125 ;
        RECT -4.340 -34.265 -4.170 -33.295 ;
        RECT -4.000 -34.085 -3.590 -33.465 ;
        RECT -3.420 -33.515 -2.920 -33.135 ;
        RECT -4.340 -34.455 -3.645 -34.265 ;
        RECT -3.420 -34.385 -3.200 -33.515 ;
        RECT -2.750 -33.685 -2.580 -32.840 ;
        RECT -1.780 -33.005 -1.610 -32.715 ;
        RECT -0.640 -32.925 -0.010 -32.675 ;
        RECT -0.180 -33.005 -0.010 -32.925 ;
        RECT 0.790 -33.005 1.030 -32.715 ;
        RECT -2.410 -33.255 -1.040 -33.005 ;
        RECT -2.410 -33.515 -2.160 -33.255 ;
        RECT -1.650 -33.685 -1.400 -33.525 ;
        RECT -2.750 -33.855 -1.400 -33.685 ;
        RECT -2.750 -33.895 -2.330 -33.855 ;
        RECT -3.020 -34.445 -2.670 -34.075 ;
        RECT -3.815 -34.785 -3.645 -34.455 ;
        RECT -2.500 -34.625 -2.330 -33.895 ;
        RECT -1.230 -34.025 -1.040 -33.255 ;
        RECT -2.160 -34.355 -1.750 -34.025 ;
        RECT -3.345 -34.825 -2.330 -34.625 ;
        RECT -1.460 -34.365 -1.040 -34.025 ;
        RECT -0.870 -33.435 -0.350 -33.125 ;
        RECT -0.180 -33.175 1.030 -33.005 ;
        RECT -0.870 -34.195 -0.700 -33.435 ;
        RECT -0.530 -34.025 -0.350 -33.615 ;
        RECT -0.180 -33.685 -0.010 -33.175 ;
        RECT 1.760 -33.325 1.930 -32.715 ;
        RECT 2.200 -33.175 2.530 -32.665 ;
        RECT 1.760 -33.345 2.080 -33.325 ;
        RECT 0.160 -33.515 2.080 -33.345 ;
        RECT -0.180 -33.855 1.720 -33.685 ;
        RECT 0.050 -34.195 0.380 -34.075 ;
        RECT -0.870 -34.365 0.380 -34.195 ;
        RECT -1.460 -34.795 -1.210 -34.365 ;
        RECT 0.550 -34.615 0.720 -33.855 ;
        RECT 1.390 -33.915 1.720 -33.855 ;
        RECT 0.910 -34.085 1.240 -34.025 ;
        RECT 0.910 -34.355 1.570 -34.085 ;
        RECT 1.890 -34.410 2.080 -33.515 ;
        RECT -0.130 -34.785 0.720 -34.615 ;
        RECT 1.760 -34.740 2.080 -34.410 ;
        RECT 2.280 -33.765 2.530 -33.175 ;
        RECT 3.175 -33.435 3.430 -32.765 ;
        RECT 3.250 -33.730 3.430 -33.435 ;
        RECT 5.875 -33.385 6.045 -32.625 ;
        RECT 5.875 -33.555 6.590 -33.385 ;
        RECT 6.760 -33.530 7.015 -32.625 ;
        RECT 3.250 -33.735 5.800 -33.730 ;
        RECT 2.280 -34.095 3.080 -33.765 ;
        RECT 2.280 -34.745 2.530 -34.095 ;
        RECT 3.250 -34.105 6.140 -33.735 ;
        RECT 6.420 -33.765 6.590 -33.555 ;
        RECT 6.420 -34.095 6.675 -33.765 ;
        RECT 3.250 -34.130 5.800 -34.105 ;
        RECT 3.250 -34.295 3.430 -34.130 ;
        RECT 6.420 -34.285 6.590 -34.095 ;
        RECT 6.845 -34.260 7.015 -33.530 ;
        RECT 37.950 -33.550 38.350 -32.050 ;
        RECT 3.175 -34.825 3.430 -34.295 ;
        RECT 5.875 -34.455 6.590 -34.285 ;
        RECT 5.875 -34.835 6.045 -34.455 ;
        RECT 6.760 -34.835 7.015 -34.260 ;
        RECT 31.495 -35.635 32.045 -35.465 ;
        RECT 31.875 -36.010 32.045 -35.635 ;
        RECT 32.225 -35.730 32.595 -35.375 ;
        RECT 32.775 -35.635 33.705 -35.465 ;
        RECT 32.775 -36.010 32.945 -35.635 ;
        RECT 31.875 -36.180 32.945 -36.010 ;
        RECT 32.235 -36.265 32.565 -36.180 ;
        RECT 31.495 -36.435 32.070 -36.350 ;
        RECT 32.800 -36.435 33.705 -36.350 ;
        RECT 31.495 -36.605 33.705 -36.435 ;
        RECT -8.535 -38.815 -8.205 -37.835 ;
        RECT 32.350 -37.950 32.550 -36.605 ;
        RECT 38.650 -37.100 39.050 -33.100 ;
        RECT 39.050 -37.550 39.350 -37.500 ;
        RECT 34.750 -37.950 39.350 -37.550 ;
        RECT -8.455 -39.030 -8.205 -38.815 ;
        RECT -0.965 -38.985 -0.585 -38.305 ;
        RECT 0.345 -38.815 0.675 -38.305 ;
        RECT 1.185 -38.815 1.585 -38.305 ;
        RECT 0.345 -38.985 1.585 -38.815 ;
        RECT -8.455 -39.200 -8.200 -39.030 ;
        RECT -8.455 -39.415 -8.205 -39.200 ;
        RECT -8.535 -40.045 -8.205 -39.415 ;
        RECT -0.965 -39.945 -0.795 -38.985 ;
        RECT -0.625 -39.325 0.680 -39.155 ;
        RECT 1.765 -39.235 2.085 -38.305 ;
        RECT 3.705 -39.065 3.875 -38.305 ;
        RECT 3.705 -39.235 4.420 -39.065 ;
        RECT 4.590 -39.210 4.845 -38.305 ;
        RECT 32.350 -38.350 35.150 -37.950 ;
        RECT 39.050 -38.000 39.350 -37.950 ;
        RECT 32.350 -38.695 32.550 -38.350 ;
        RECT 32.315 -39.025 32.565 -38.695 ;
        RECT 39.550 -38.700 39.950 -33.100 ;
        RECT 40.450 -37.100 40.850 -32.050 ;
        RECT 40.150 -38.000 40.450 -37.500 ;
        RECT 43.450 -38.700 43.850 -33.250 ;
        RECT 44.350 -35.250 44.750 -31.050 ;
        RECT 45.250 -35.250 45.650 -33.250 ;
        RECT 47.300 -35.250 47.700 -33.250 ;
        RECT 48.200 -35.250 48.600 -31.050 ;
        RECT 51.800 -31.550 52.200 -31.050 ;
        RECT 51.800 -32.050 52.900 -31.550 ;
        RECT 44.050 -36.150 45.050 -35.650 ;
        RECT 48.000 -36.150 48.850 -35.650 ;
        RECT 39.550 -39.100 43.850 -38.700 ;
        RECT -0.625 -39.775 -0.380 -39.325 ;
        RECT -0.210 -39.695 0.340 -39.495 ;
        RECT 0.510 -39.525 0.680 -39.325 ;
        RECT 1.455 -39.380 2.085 -39.235 ;
        RECT 1.455 -39.430 3.300 -39.380 ;
        RECT 3.615 -39.430 3.970 -39.415 ;
        RECT 0.510 -39.695 0.885 -39.525 ;
        RECT 1.055 -39.945 1.285 -39.445 ;
        RECT -0.965 -40.115 1.285 -39.945 ;
        RECT 1.455 -39.630 3.970 -39.430 ;
        RECT -0.415 -40.435 -0.245 -40.115 ;
        RECT 1.455 -40.285 1.625 -39.630 ;
        RECT 3.615 -39.785 3.970 -39.630 ;
        RECT 4.250 -39.445 4.420 -39.235 ;
        RECT 4.250 -39.775 4.505 -39.445 ;
        RECT 4.250 -39.965 4.420 -39.775 ;
        RECT 4.675 -39.940 4.845 -39.210 ;
        RECT 31.495 -39.195 32.125 -39.115 ;
        RECT 32.725 -39.195 33.705 -39.115 ;
        RECT 6.300 -39.750 11.850 -39.350 ;
        RECT 31.495 -39.445 33.705 -39.195 ;
        RECT 44.350 -39.500 44.750 -36.150 ;
        RECT 49.100 -38.350 49.500 -33.250 ;
        RECT 51.800 -33.700 52.200 -32.050 ;
        RECT 52.500 -37.150 52.900 -32.050 ;
        RECT 52.900 -38.050 53.200 -37.550 ;
        RECT 53.400 -38.350 53.800 -33.150 ;
        RECT 54.300 -37.150 54.700 -33.150 ;
        RECT 54.000 -38.050 54.300 -37.550 ;
        RECT 55.900 -38.350 56.400 -27.900 ;
        RECT 70.400 -27.875 71.425 -27.625 ;
        RECT 65.685 -29.605 66.015 -28.795 ;
        RECT 65.685 -29.775 66.400 -29.605 ;
        RECT 65.680 -29.950 66.060 -29.945 ;
        RECT 64.100 -30.150 66.060 -29.950 ;
        RECT 64.100 -32.300 64.400 -30.150 ;
        RECT 65.680 -30.185 66.060 -30.150 ;
        RECT 66.230 -30.015 66.400 -29.775 ;
        RECT 66.605 -29.645 66.775 -28.795 ;
        RECT 67.445 -29.645 67.615 -28.795 ;
        RECT 70.400 -29.150 70.650 -27.875 ;
        RECT 66.605 -29.815 67.615 -29.645 ;
        RECT 67.120 -29.950 67.615 -29.815 ;
        RECT 68.350 -29.400 70.650 -29.150 ;
        RECT 71.165 -29.295 71.335 -28.795 ;
        RECT 68.350 -29.950 68.625 -29.400 ;
        RECT 71.165 -29.465 71.830 -29.295 ;
        RECT 66.230 -30.185 66.730 -30.015 ;
        RECT 66.230 -30.355 66.400 -30.185 ;
        RECT 67.120 -30.200 68.625 -29.950 ;
        RECT 67.120 -30.355 67.615 -30.200 ;
        RECT 71.080 -30.285 71.430 -29.635 ;
        RECT 65.765 -30.525 66.400 -30.355 ;
        RECT 66.605 -30.525 67.615 -30.355 ;
        RECT 71.600 -30.455 71.830 -29.465 ;
        RECT 65.765 -31.005 65.935 -30.525 ;
        RECT 66.605 -31.005 66.775 -30.525 ;
        RECT 67.445 -31.005 67.615 -30.525 ;
        RECT 71.165 -30.625 71.830 -30.455 ;
        RECT 71.165 -30.915 71.335 -30.625 ;
        RECT 72.005 -30.915 72.190 -28.795 ;
        RECT 72.865 -29.220 73.115 -28.795 ;
        RECT 73.325 -29.070 74.430 -28.900 ;
        RECT 72.810 -29.350 73.115 -29.220 ;
        RECT 72.360 -30.545 72.640 -29.595 ;
        RECT 72.810 -30.455 72.980 -29.350 ;
        RECT 73.150 -30.135 73.390 -29.540 ;
        RECT 73.560 -29.605 74.090 -29.240 ;
        RECT 73.560 -30.305 73.730 -29.605 ;
        RECT 74.260 -29.685 74.430 -29.070 ;
        RECT 74.940 -29.125 75.190 -28.795 ;
        RECT 75.415 -29.095 76.300 -28.925 ;
        RECT 74.260 -29.775 74.770 -29.685 ;
        RECT 72.810 -30.585 73.035 -30.455 ;
        RECT 73.205 -30.525 73.730 -30.305 ;
        RECT 73.900 -29.945 74.770 -29.775 ;
        RECT 72.865 -30.725 73.035 -30.585 ;
        RECT 73.900 -30.725 74.070 -29.945 ;
        RECT 74.600 -30.015 74.770 -29.945 ;
        RECT 74.280 -30.195 74.480 -30.165 ;
        RECT 74.940 -30.195 75.110 -29.125 ;
        RECT 75.280 -30.015 75.470 -29.295 ;
        RECT 74.280 -30.495 75.110 -30.195 ;
        RECT 75.640 -30.225 75.960 -29.265 ;
        RECT 72.865 -30.895 73.200 -30.725 ;
        RECT 73.395 -30.895 74.070 -30.725 ;
        RECT 74.940 -30.725 75.110 -30.495 ;
        RECT 75.495 -30.555 75.960 -30.225 ;
        RECT 76.130 -29.935 76.300 -29.095 ;
        RECT 77.030 -29.355 77.370 -28.795 ;
        RECT 76.470 -29.730 77.370 -29.355 ;
        RECT 77.180 -29.935 77.370 -29.730 ;
        RECT 77.880 -29.685 78.210 -28.840 ;
        RECT 78.895 -29.545 79.225 -28.815 ;
        RECT 77.880 -29.765 78.290 -29.685 ;
        RECT 78.055 -29.815 78.290 -29.765 ;
        RECT 76.130 -30.265 77.010 -29.935 ;
        RECT 77.180 -30.265 77.930 -29.935 ;
        RECT 76.130 -30.725 76.300 -30.265 ;
        RECT 77.180 -30.435 77.380 -30.265 ;
        RECT 78.100 -30.395 78.290 -29.815 ;
        RECT 78.045 -30.435 78.290 -30.395 ;
        RECT 74.940 -30.895 75.345 -30.725 ;
        RECT 75.515 -30.895 76.300 -30.725 ;
        RECT 77.050 -30.960 77.380 -30.435 ;
        RECT 77.890 -30.520 78.290 -30.435 ;
        RECT 78.955 -29.935 79.225 -29.545 ;
        RECT 79.800 -29.765 80.135 -28.795 ;
        RECT 78.955 -30.265 79.750 -29.935 ;
        RECT 79.920 -29.950 80.135 -29.765 ;
        RECT 79.920 -30.150 82.100 -29.950 ;
        RECT 77.890 -30.955 78.220 -30.520 ;
        RECT 78.955 -30.645 79.155 -30.265 ;
        RECT 79.920 -30.375 80.135 -30.150 ;
        RECT 80.750 -30.300 82.100 -30.150 ;
        RECT 78.895 -30.915 79.155 -30.645 ;
        RECT 79.880 -30.995 80.135 -30.375 ;
        RECT 80.900 -30.900 81.400 -30.500 ;
        RECT 81.700 -32.300 82.100 -30.300 ;
        RECT 64.100 -32.700 82.100 -32.300 ;
        RECT 68.355 -37.095 68.685 -36.295 ;
        RECT 69.195 -37.075 69.525 -36.295 ;
        RECT 72.565 -36.795 72.735 -36.295 ;
        RECT 72.565 -36.965 73.230 -36.795 ;
        RECT 69.195 -37.095 69.960 -37.075 ;
        RECT 68.355 -37.150 69.960 -37.095 ;
        RECT 72.480 -37.150 72.830 -37.135 ;
        RECT 68.355 -37.265 72.830 -37.150 ;
        RECT 67.895 -37.685 69.525 -37.435 ;
        RECT 69.695 -37.550 72.830 -37.265 ;
        RECT 69.695 -37.855 69.960 -37.550 ;
        RECT 72.480 -37.785 72.830 -37.550 ;
        RECT 49.100 -38.850 56.400 -38.350 ;
        RECT 68.355 -38.035 69.960 -37.855 ;
        RECT 73.000 -37.955 73.230 -36.965 ;
        RECT 68.355 -38.505 68.685 -38.035 ;
        RECT 69.195 -38.505 69.525 -38.035 ;
        RECT 71.000 -38.450 71.550 -38.000 ;
        RECT 72.565 -38.125 73.230 -37.955 ;
        RECT 72.565 -38.415 72.735 -38.125 ;
        RECT 73.405 -38.415 73.590 -36.295 ;
        RECT 74.265 -36.720 74.515 -36.295 ;
        RECT 74.725 -36.570 75.830 -36.400 ;
        RECT 74.210 -36.850 74.515 -36.720 ;
        RECT 73.760 -38.045 74.040 -37.095 ;
        RECT 74.210 -37.955 74.380 -36.850 ;
        RECT 74.550 -37.635 74.790 -37.040 ;
        RECT 74.960 -37.105 75.490 -36.740 ;
        RECT 74.960 -37.805 75.130 -37.105 ;
        RECT 75.660 -37.185 75.830 -36.570 ;
        RECT 76.340 -36.625 76.590 -36.295 ;
        RECT 76.815 -36.595 77.700 -36.425 ;
        RECT 75.660 -37.275 76.170 -37.185 ;
        RECT 74.210 -38.085 74.435 -37.955 ;
        RECT 74.605 -38.025 75.130 -37.805 ;
        RECT 75.300 -37.445 76.170 -37.275 ;
        RECT 74.265 -38.225 74.435 -38.085 ;
        RECT 75.300 -38.225 75.470 -37.445 ;
        RECT 76.000 -37.515 76.170 -37.445 ;
        RECT 75.680 -37.695 75.880 -37.665 ;
        RECT 76.340 -37.695 76.510 -36.625 ;
        RECT 76.680 -37.515 76.870 -36.795 ;
        RECT 75.680 -37.995 76.510 -37.695 ;
        RECT 77.040 -37.725 77.360 -36.765 ;
        RECT 74.265 -38.395 74.600 -38.225 ;
        RECT 74.795 -38.395 75.470 -38.225 ;
        RECT 76.340 -38.225 76.510 -37.995 ;
        RECT 76.895 -38.055 77.360 -37.725 ;
        RECT 77.530 -37.435 77.700 -36.595 ;
        RECT 78.425 -36.855 78.765 -36.295 ;
        RECT 77.870 -37.230 78.765 -36.855 ;
        RECT 78.575 -37.435 78.765 -37.230 ;
        RECT 79.275 -37.185 79.605 -36.340 ;
        RECT 79.275 -37.265 79.665 -37.185 ;
        RECT 79.450 -37.315 79.665 -37.265 ;
        RECT 77.530 -37.765 78.405 -37.435 ;
        RECT 78.575 -37.765 79.325 -37.435 ;
        RECT 77.530 -38.225 77.700 -37.765 ;
        RECT 78.575 -37.935 78.775 -37.765 ;
        RECT 79.495 -37.895 79.665 -37.315 ;
        RECT 79.440 -37.935 79.665 -37.895 ;
        RECT 76.340 -38.395 76.745 -38.225 ;
        RECT 76.915 -38.395 77.700 -38.225 ;
        RECT 71.175 -39.325 71.425 -38.450 ;
        RECT 78.445 -38.460 78.775 -37.935 ;
        RECT 79.285 -38.020 79.665 -37.935 ;
        RECT 79.285 -38.455 79.615 -38.020 ;
        RECT 0.670 -40.455 1.625 -40.285 ;
        RECT 3.705 -40.135 4.420 -39.965 ;
        RECT 3.705 -40.515 3.875 -40.135 ;
        RECT 4.590 -40.515 4.845 -39.940 ;
        RECT 34.750 -40.000 54.700 -39.500 ;
        RECT 70.400 -39.575 71.425 -39.325 ;
        RECT 34.750 -40.600 35.250 -40.000 ;
        RECT 32.600 -41.100 35.250 -40.600 ;
        RECT 65.685 -41.305 66.015 -40.495 ;
        RECT 65.685 -41.475 66.400 -41.305 ;
        RECT 65.680 -41.650 66.060 -41.645 ;
        RECT 64.100 -41.850 66.060 -41.650 ;
        RECT 40.830 -42.820 42.990 -42.470 ;
        RECT -7.675 -43.625 -7.345 -42.995 ;
        RECT -5.270 -43.535 -5.015 -43.005 ;
        RECT -7.675 -44.225 -7.425 -43.625 ;
        RECT -7.255 -43.820 -6.925 -43.815 ;
        RECT -5.270 -43.820 -5.090 -43.535 ;
        RECT -4.370 -43.735 -4.120 -43.085 ;
        RECT -7.255 -44.060 -5.090 -43.820 ;
        RECT -7.255 -44.065 -6.925 -44.060 ;
        RECT -7.675 -45.205 -7.345 -44.225 ;
        RECT -5.270 -44.395 -5.090 -44.060 ;
        RECT -4.920 -44.065 -4.120 -43.735 ;
        RECT -5.270 -45.065 -5.015 -44.395 ;
        RECT -4.370 -44.655 -4.120 -44.065 ;
        RECT -3.920 -43.420 -3.600 -43.090 ;
        RECT -2.560 -43.215 -1.710 -43.045 ;
        RECT -3.920 -44.315 -3.730 -43.420 ;
        RECT -3.410 -43.745 -2.750 -43.475 ;
        RECT -3.080 -43.805 -2.750 -43.745 ;
        RECT -3.560 -43.975 -3.230 -43.915 ;
        RECT -2.560 -43.975 -2.390 -43.215 ;
        RECT -0.630 -43.465 -0.380 -43.035 ;
        RECT -2.220 -43.635 -0.970 -43.465 ;
        RECT -2.220 -43.755 -1.890 -43.635 ;
        RECT -3.560 -44.145 -1.660 -43.975 ;
        RECT -3.920 -44.485 -2.000 -44.315 ;
        RECT -3.920 -44.505 -3.600 -44.485 ;
        RECT -4.370 -45.165 -4.040 -44.655 ;
        RECT -3.770 -45.115 -3.600 -44.505 ;
        RECT -1.830 -44.655 -1.660 -44.145 ;
        RECT -1.490 -44.215 -1.310 -43.805 ;
        RECT -1.140 -44.395 -0.970 -43.635 ;
        RECT -2.870 -44.825 -1.660 -44.655 ;
        RECT -1.490 -44.705 -0.970 -44.395 ;
        RECT -0.800 -43.805 -0.380 -43.465 ;
        RECT 0.490 -43.205 1.505 -43.005 ;
        RECT -0.090 -43.805 0.320 -43.475 ;
        RECT -0.800 -44.575 -0.610 -43.805 ;
        RECT 0.490 -43.935 0.660 -43.205 ;
        RECT 1.805 -43.375 1.975 -43.045 ;
        RECT 0.830 -43.755 1.180 -43.385 ;
        RECT 0.490 -43.975 0.910 -43.935 ;
        RECT -0.440 -44.145 0.910 -43.975 ;
        RECT -0.440 -44.305 -0.190 -44.145 ;
        RECT 0.320 -44.575 0.570 -44.315 ;
        RECT -0.800 -44.825 0.570 -44.575 ;
        RECT -2.870 -45.115 -2.630 -44.825 ;
        RECT -1.830 -44.905 -1.660 -44.825 ;
        RECT -1.830 -45.155 -1.200 -44.905 ;
        RECT -0.230 -45.115 -0.060 -44.825 ;
        RECT 0.740 -44.990 0.910 -44.145 ;
        RECT 1.360 -44.315 1.580 -43.445 ;
        RECT 1.805 -43.565 2.500 -43.375 ;
        RECT 1.080 -44.695 1.580 -44.315 ;
        RECT 1.750 -44.365 2.160 -43.745 ;
        RECT 2.330 -44.535 2.500 -43.565 ;
        RECT 1.805 -44.705 2.500 -44.535 ;
        RECT 0.740 -45.160 1.570 -44.990 ;
        RECT 1.805 -45.205 1.975 -44.705 ;
        RECT 2.690 -45.205 2.915 -43.085 ;
        RECT 3.585 -43.375 3.755 -43.085 ;
        RECT 3.090 -43.545 3.755 -43.375 ;
        RECT 3.090 -44.535 3.320 -43.545 ;
        RECT 6.385 -43.570 6.640 -42.995 ;
        RECT 7.355 -43.375 7.525 -42.995 ;
        RECT 6.810 -43.545 7.525 -43.375 ;
        RECT 3.490 -43.730 3.840 -43.715 ;
        RECT 3.490 -44.080 5.400 -43.730 ;
        RECT 3.490 -44.365 3.840 -44.080 ;
        RECT 6.385 -44.300 6.555 -43.570 ;
        RECT 6.810 -43.735 6.980 -43.545 ;
        RECT 19.250 -43.650 19.750 -43.150 ;
        RECT 7.900 -43.720 19.750 -43.650 ;
        RECT 6.725 -44.065 6.980 -43.735 ;
        RECT 6.810 -44.275 6.980 -44.065 ;
        RECT 7.260 -44.100 19.750 -43.720 ;
        RECT 7.900 -44.150 19.750 -44.100 ;
        RECT 64.100 -44.000 64.400 -41.850 ;
        RECT 65.680 -41.885 66.060 -41.850 ;
        RECT 66.230 -41.715 66.400 -41.475 ;
        RECT 66.605 -41.345 66.775 -40.495 ;
        RECT 67.445 -41.345 67.615 -40.495 ;
        RECT 70.400 -40.850 70.650 -39.575 ;
        RECT 81.400 -39.850 85.850 -39.350 ;
        RECT 81.400 -40.250 81.900 -39.850 ;
        RECT 66.605 -41.515 67.615 -41.345 ;
        RECT 67.120 -41.650 67.615 -41.515 ;
        RECT 68.350 -41.100 70.650 -40.850 ;
        RECT 71.165 -40.995 71.335 -40.495 ;
        RECT 68.350 -41.650 68.625 -41.100 ;
        RECT 71.165 -41.165 71.830 -40.995 ;
        RECT 66.230 -41.885 66.730 -41.715 ;
        RECT 66.230 -42.055 66.400 -41.885 ;
        RECT 67.120 -41.900 68.625 -41.650 ;
        RECT 67.120 -42.055 67.615 -41.900 ;
        RECT 71.080 -41.985 71.430 -41.335 ;
        RECT 65.765 -42.225 66.400 -42.055 ;
        RECT 66.605 -42.225 67.615 -42.055 ;
        RECT 71.600 -42.155 71.830 -41.165 ;
        RECT 65.765 -42.705 65.935 -42.225 ;
        RECT 66.605 -42.705 66.775 -42.225 ;
        RECT 67.445 -42.705 67.615 -42.225 ;
        RECT 71.165 -42.325 71.830 -42.155 ;
        RECT 71.165 -42.615 71.335 -42.325 ;
        RECT 72.005 -42.615 72.190 -40.495 ;
        RECT 72.865 -40.920 73.115 -40.495 ;
        RECT 73.325 -40.770 74.430 -40.600 ;
        RECT 72.810 -41.050 73.115 -40.920 ;
        RECT 72.360 -42.245 72.640 -41.295 ;
        RECT 72.810 -42.155 72.980 -41.050 ;
        RECT 73.150 -41.835 73.390 -41.240 ;
        RECT 73.560 -41.305 74.090 -40.940 ;
        RECT 73.560 -42.005 73.730 -41.305 ;
        RECT 74.260 -41.385 74.430 -40.770 ;
        RECT 74.940 -40.825 75.190 -40.495 ;
        RECT 75.415 -40.795 76.300 -40.625 ;
        RECT 74.260 -41.475 74.770 -41.385 ;
        RECT 72.810 -42.285 73.035 -42.155 ;
        RECT 73.205 -42.225 73.730 -42.005 ;
        RECT 73.900 -41.645 74.770 -41.475 ;
        RECT 72.865 -42.425 73.035 -42.285 ;
        RECT 73.900 -42.425 74.070 -41.645 ;
        RECT 74.600 -41.715 74.770 -41.645 ;
        RECT 74.280 -41.895 74.480 -41.865 ;
        RECT 74.940 -41.895 75.110 -40.825 ;
        RECT 75.280 -41.715 75.470 -40.995 ;
        RECT 74.280 -42.195 75.110 -41.895 ;
        RECT 75.640 -41.925 75.960 -40.965 ;
        RECT 72.865 -42.595 73.200 -42.425 ;
        RECT 73.395 -42.595 74.070 -42.425 ;
        RECT 74.940 -42.425 75.110 -42.195 ;
        RECT 75.495 -42.255 75.960 -41.925 ;
        RECT 76.130 -41.635 76.300 -40.795 ;
        RECT 77.030 -41.055 77.370 -40.495 ;
        RECT 76.470 -41.430 77.370 -41.055 ;
        RECT 77.180 -41.635 77.370 -41.430 ;
        RECT 77.880 -41.385 78.210 -40.540 ;
        RECT 78.895 -41.245 79.225 -40.515 ;
        RECT 77.880 -41.465 78.290 -41.385 ;
        RECT 78.055 -41.515 78.290 -41.465 ;
        RECT 76.130 -41.965 77.010 -41.635 ;
        RECT 77.180 -41.965 77.930 -41.635 ;
        RECT 76.130 -42.425 76.300 -41.965 ;
        RECT 77.180 -42.135 77.380 -41.965 ;
        RECT 78.100 -42.095 78.290 -41.515 ;
        RECT 78.045 -42.135 78.290 -42.095 ;
        RECT 74.940 -42.595 75.345 -42.425 ;
        RECT 75.515 -42.595 76.300 -42.425 ;
        RECT 77.050 -42.660 77.380 -42.135 ;
        RECT 77.890 -42.220 78.290 -42.135 ;
        RECT 78.955 -41.635 79.225 -41.245 ;
        RECT 79.800 -41.465 80.135 -40.495 ;
        RECT 78.955 -41.965 79.750 -41.635 ;
        RECT 79.920 -41.650 80.135 -41.465 ;
        RECT 79.920 -41.850 82.100 -41.650 ;
        RECT 77.890 -42.655 78.220 -42.220 ;
        RECT 78.955 -42.345 79.155 -41.965 ;
        RECT 79.920 -42.075 80.135 -41.850 ;
        RECT 80.750 -42.000 82.100 -41.850 ;
        RECT 78.895 -42.615 79.155 -42.345 ;
        RECT 79.880 -42.695 80.135 -42.075 ;
        RECT 80.900 -42.600 81.400 -42.200 ;
        RECT 81.700 -44.000 82.100 -42.000 ;
        RECT 3.090 -44.705 3.755 -44.535 ;
        RECT 3.585 -45.205 3.755 -44.705 ;
        RECT 6.385 -45.205 6.640 -44.300 ;
        RECT 6.810 -44.445 7.525 -44.275 ;
        RECT 64.100 -44.400 82.100 -44.000 ;
        RECT 7.355 -45.205 7.525 -44.445 ;
        RECT 85.350 -50.100 85.850 -39.850 ;
        RECT 85.000 -50.500 85.850 -50.100 ;
      LAYER met1 ;
        RECT -2.150 37.450 -1.750 37.950 ;
        RECT 12.800 37.450 13.200 37.950 ;
        RECT 27.850 37.450 28.250 37.950 ;
        RECT 42.800 37.450 43.200 37.950 ;
        RECT 57.850 37.450 58.250 37.950 ;
        RECT 72.800 37.450 73.200 37.950 ;
        RECT -10.100 36.950 -3.100 37.450 ;
        RECT -10.100 10.100 -9.600 36.950 ;
        RECT -3.600 33.850 -3.100 36.950 ;
        RECT -2.150 36.950 26.900 37.450 ;
        RECT -2.150 36.550 -1.750 36.950 ;
        RECT 5.200 33.850 5.700 36.950 ;
        RECT 12.800 36.550 13.200 36.950 ;
        RECT 7.350 35.900 7.750 36.250 ;
        RECT 18.250 35.900 18.650 36.250 ;
        RECT 7.350 35.400 18.650 35.900 ;
        RECT 7.350 35.050 7.750 35.400 ;
        RECT 10.050 33.850 10.550 35.400 ;
        RECT 18.250 35.050 18.650 35.400 ;
        RECT 26.400 33.850 26.900 36.950 ;
        RECT 27.850 36.950 56.900 37.450 ;
        RECT 27.850 36.550 28.250 36.950 ;
        RECT 35.200 33.850 35.700 36.950 ;
        RECT 42.800 36.550 43.200 36.950 ;
        RECT 37.350 35.900 37.750 36.250 ;
        RECT 48.250 35.900 48.650 36.250 ;
        RECT 37.350 35.400 48.650 35.900 ;
        RECT 37.350 35.050 37.750 35.400 ;
        RECT 40.050 33.850 40.550 35.400 ;
        RECT 48.250 35.050 48.650 35.400 ;
        RECT 56.400 33.850 56.900 36.950 ;
        RECT 57.850 36.950 87.800 37.450 ;
        RECT 57.850 36.550 58.250 36.950 ;
        RECT 65.200 33.850 65.700 36.950 ;
        RECT 72.800 36.550 73.200 36.950 ;
        RECT 67.350 35.900 67.750 36.250 ;
        RECT 78.250 35.900 78.650 36.250 ;
        RECT 67.350 35.400 78.650 35.900 ;
        RECT 67.350 35.050 67.750 35.400 ;
        RECT 70.050 33.850 70.550 35.400 ;
        RECT 78.250 35.050 78.650 35.400 ;
        RECT -5.000 33.200 -0.100 33.850 ;
        RECT 4.850 33.200 6.050 33.850 ;
        RECT 9.700 33.200 10.900 33.850 ;
        RECT 15.400 33.750 20.300 33.850 ;
        RECT 14.550 33.250 20.300 33.750 ;
        RECT 14.550 31.100 15.050 33.250 ;
        RECT 15.400 33.200 20.300 33.250 ;
        RECT 25.000 33.200 29.900 33.850 ;
        RECT 34.850 33.200 36.050 33.850 ;
        RECT 39.700 33.200 40.900 33.850 ;
        RECT 45.400 33.750 50.300 33.850 ;
        RECT 44.550 33.250 50.300 33.750 ;
        RECT -8.600 30.600 15.050 31.100 ;
        RECT 18.250 31.100 18.650 31.400 ;
        RECT 44.550 31.100 45.050 33.250 ;
        RECT 45.400 33.200 50.300 33.250 ;
        RECT 55.000 33.200 59.900 33.850 ;
        RECT 64.850 33.200 66.050 33.850 ;
        RECT 69.700 33.200 70.900 33.850 ;
        RECT 75.400 33.750 80.300 33.850 ;
        RECT 74.550 33.250 80.300 33.750 ;
        RECT 18.250 30.600 45.050 31.100 ;
        RECT 48.250 31.100 48.650 31.400 ;
        RECT 74.550 31.100 75.050 33.250 ;
        RECT 75.400 33.200 80.300 33.250 ;
        RECT 48.250 30.600 75.050 31.100 ;
        RECT 78.250 31.100 78.650 31.400 ;
        RECT 78.250 30.600 84.900 31.100 ;
        RECT -8.600 16.450 -8.100 30.600 ;
        RECT 18.250 30.200 18.650 30.600 ;
        RECT 48.250 30.200 48.650 30.600 ;
        RECT 78.250 30.200 78.650 30.600 ;
        RECT 24.970 24.250 27.075 24.630 ;
        RECT 24.970 22.700 27.075 23.080 ;
        RECT 17.300 19.200 17.750 19.300 ;
        RECT 14.350 18.900 17.750 19.200 ;
        RECT 14.350 16.450 14.850 18.900 ;
        RECT 17.300 18.850 17.750 18.900 ;
        RECT 27.150 16.450 27.550 16.850 ;
        RECT 57.150 16.450 57.550 16.850 ;
        RECT 83.900 16.450 84.900 30.600 ;
        RECT -8.600 15.950 27.550 16.450 ;
        RECT 27.150 15.650 27.550 15.950 ;
        RECT 30.750 15.950 57.550 16.450 ;
        RECT 25.500 13.800 30.400 13.850 ;
        RECT 30.750 13.800 31.250 15.950 ;
        RECT 57.150 15.650 57.550 15.950 ;
        RECT 60.750 15.950 84.900 16.450 ;
        RECT 25.500 13.300 31.250 13.800 ;
        RECT 25.500 13.200 30.400 13.300 ;
        RECT 34.900 13.200 36.100 13.850 ;
        RECT 39.750 13.200 40.950 13.850 ;
        RECT 45.900 13.200 50.800 13.850 ;
        RECT 55.500 13.800 60.400 13.850 ;
        RECT 60.750 13.800 61.250 15.950 ;
        RECT 55.500 13.300 61.250 13.800 ;
        RECT 55.500 13.200 60.400 13.300 ;
        RECT 64.900 13.200 66.100 13.850 ;
        RECT 69.750 13.200 70.950 13.850 ;
        RECT 75.900 13.200 80.800 13.850 ;
        RECT 27.150 11.650 27.550 12.000 ;
        RECT 35.250 11.650 35.750 13.200 ;
        RECT 38.050 11.650 38.450 12.000 ;
        RECT 27.150 11.150 38.450 11.650 ;
        RECT 27.150 10.800 27.550 11.150 ;
        RECT 38.050 10.800 38.450 11.150 ;
        RECT 32.600 10.100 33.000 10.500 ;
        RECT 40.100 10.100 40.600 13.200 ;
        RECT 47.550 10.100 47.950 10.500 ;
        RECT -10.100 9.600 47.950 10.100 ;
        RECT 48.900 10.100 49.400 13.200 ;
        RECT 57.150 11.650 57.550 12.000 ;
        RECT 65.250 11.650 65.750 13.200 ;
        RECT 68.050 11.650 68.450 12.000 ;
        RECT 57.150 11.150 68.450 11.650 ;
        RECT 57.150 10.800 57.550 11.150 ;
        RECT 68.050 10.800 68.450 11.150 ;
        RECT 62.600 10.100 63.000 10.500 ;
        RECT 70.100 10.100 70.600 13.200 ;
        RECT 77.550 10.100 77.950 10.500 ;
        RECT 48.900 9.600 77.950 10.100 ;
        RECT 78.900 10.100 79.400 13.200 ;
        RECT 86.800 10.100 87.800 36.950 ;
        RECT 78.900 9.600 87.800 10.100 ;
        RECT -10.100 -2.050 -9.600 9.600 ;
        RECT 32.600 9.100 33.000 9.600 ;
        RECT 47.550 9.100 47.950 9.600 ;
        RECT 62.600 9.100 63.000 9.600 ;
        RECT 77.550 9.100 77.950 9.600 ;
        RECT 79.800 3.550 86.800 3.950 ;
        RECT 34.600 2.200 35.000 2.700 ;
        RECT 39.300 2.100 39.700 2.600 ;
        RECT 42.400 2.100 42.800 2.600 ;
        RECT 45.500 2.200 45.900 2.700 ;
        RECT 50.200 2.200 50.600 2.700 ;
        RECT 54.900 2.100 55.300 2.600 ;
        RECT 58.000 2.100 58.400 2.600 ;
        RECT 61.100 2.200 61.500 2.700 ;
        RECT 65.800 2.200 66.200 2.700 ;
        RECT 70.500 2.100 70.900 2.600 ;
        RECT 73.600 2.100 74.000 2.600 ;
        RECT 76.700 2.200 77.100 2.700 ;
        RECT 36.900 1.650 37.300 1.850 ;
        RECT 44.700 1.650 45.100 1.850 ;
        RECT 36.900 1.450 45.100 1.650 ;
        RECT 52.500 1.650 52.900 1.850 ;
        RECT 60.300 1.650 60.700 1.850 ;
        RECT 52.500 1.450 60.700 1.650 ;
        RECT 68.100 1.650 68.500 1.850 ;
        RECT 75.900 1.650 76.300 1.850 ;
        RECT 68.100 1.450 76.300 1.650 ;
        RECT 31.900 1.050 36.350 1.450 ;
        RECT 36.900 1.250 51.950 1.450 ;
        RECT 36.900 1.050 37.300 1.250 ;
        RECT -5.220 -1.500 -4.930 -1.455 ;
        RECT -3.360 -1.500 -3.070 -1.455 ;
        RECT -0.580 -1.500 -0.290 -1.455 ;
        RECT -5.220 -1.640 -0.290 -1.500 ;
        RECT -5.220 -1.685 -4.930 -1.640 ;
        RECT -3.360 -1.685 -3.070 -1.640 ;
        RECT -0.580 -1.685 -0.290 -1.640 ;
        RECT 6.750 -1.680 9.050 -1.330 ;
        RECT -10.100 -2.450 -9.300 -2.050 ;
        RECT -6.750 -2.330 -3.600 -1.930 ;
        RECT -0.580 -2.180 -0.290 -2.135 ;
        RECT -2.825 -2.320 -0.290 -2.180 ;
        RECT -8.050 -7.280 -7.600 -7.230 ;
        RECT -8.450 -7.630 -7.600 -7.280 ;
        RECT -8.050 -7.680 -7.600 -7.630 ;
        RECT -6.750 -9.180 -6.400 -2.330 ;
        RECT -2.825 -2.475 -2.610 -2.320 ;
        RECT -0.580 -2.365 -0.290 -2.320 ;
        RECT -4.760 -2.520 -4.470 -2.475 ;
        RECT -2.900 -2.520 -2.610 -2.475 ;
        RECT -1.980 -2.480 -1.690 -2.475 ;
        RECT -4.760 -2.660 -2.610 -2.520 ;
        RECT -4.760 -2.705 -4.470 -2.660 ;
        RECT -2.900 -2.705 -2.610 -2.660 ;
        RECT -2.050 -2.520 -1.550 -2.480 ;
        RECT 1.280 -2.520 1.570 -2.475 ;
        RECT -2.050 -2.660 1.570 -2.520 ;
        RECT -2.050 -2.930 -1.550 -2.660 ;
        RECT 1.280 -2.705 1.570 -2.660 ;
        RECT 4.700 -4.930 5.050 -2.080 ;
        RECT -2.650 -5.280 5.050 -4.930 ;
        RECT -2.650 -6.930 -2.300 -5.280 ;
        RECT -2.650 -7.280 0.250 -6.930 ;
        RECT -0.700 -8.130 -0.350 -7.780 ;
        RECT -0.100 -7.830 0.250 -7.280 ;
        RECT 4.550 -7.700 4.850 -7.030 ;
        RECT -0.200 -8.080 0.350 -7.830 ;
        RECT 4.550 -8.090 6.450 -7.700 ;
        RECT 4.850 -8.100 6.450 -8.090 ;
        RECT -9.400 -9.480 -6.400 -9.180 ;
        RECT -2.650 -8.480 -0.350 -8.130 ;
        RECT -9.400 -11.630 -9.050 -9.480 ;
        RECT -2.650 -10.180 -2.300 -8.480 ;
        RECT 8.700 -9.980 9.050 -1.680 ;
        RECT 29.750 -8.100 30.550 -7.700 ;
        RECT -6.400 -10.530 -2.300 -10.180 ;
        RECT 4.350 -10.330 9.050 -9.980 ;
        RECT -6.400 -11.580 -6.050 -10.530 ;
        RECT -9.400 -11.980 -7.350 -11.630 ;
        RECT -6.400 -11.980 -4.950 -11.580 ;
        RECT -3.410 -11.870 -3.120 -11.825 ;
        RECT -0.150 -11.870 0.350 -11.530 ;
        RECT -3.410 -12.010 0.350 -11.870 ;
        RECT -3.410 -12.055 -3.120 -12.010 ;
        RECT -0.150 -12.030 0.350 -12.010 ;
        RECT 0.770 -11.870 1.060 -11.825 ;
        RECT 2.630 -11.870 2.920 -11.825 ;
        RECT 0.770 -12.010 2.920 -11.870 ;
        RECT -0.150 -12.055 0.140 -12.030 ;
        RECT 0.770 -12.055 1.060 -12.010 ;
        RECT 2.630 -12.055 2.920 -12.010 ;
        RECT -1.550 -12.210 -1.260 -12.165 ;
        RECT 0.770 -12.210 0.985 -12.055 ;
        RECT -1.550 -12.350 0.985 -12.210 ;
        RECT -1.550 -12.395 -1.260 -12.350 ;
        RECT 1.750 -12.380 2.150 -12.180 ;
        RECT 4.350 -12.380 4.700 -10.330 ;
        RECT 1.750 -12.680 4.700 -12.380 ;
        RECT 5.050 -12.430 6.700 -12.080 ;
        RECT 1.750 -12.730 2.950 -12.680 ;
        RECT 3.550 -12.730 4.700 -12.680 ;
        RECT -1.550 -12.890 -1.260 -12.845 ;
        RECT 1.230 -12.890 1.520 -12.845 ;
        RECT 3.090 -12.890 3.380 -12.845 ;
        RECT -1.550 -13.030 3.380 -12.890 ;
        RECT -1.550 -13.075 -1.260 -13.030 ;
        RECT 1.230 -13.075 1.520 -13.030 ;
        RECT 3.090 -13.075 3.380 -13.030 ;
        RECT 6.350 -13.230 6.700 -12.430 ;
        RECT 18.750 -12.500 19.750 -12.000 ;
        RECT -6.380 -25.010 -6.080 -24.160 ;
        RECT 8.800 -24.400 9.200 -24.250 ;
        RECT 10.400 -24.400 12.100 -24.350 ;
        RECT -3.040 -24.520 -2.750 -24.475 ;
        RECT -0.940 -24.520 -0.650 -24.475 ;
        RECT 0.630 -24.520 0.920 -24.475 ;
        RECT -3.040 -24.660 0.920 -24.520 ;
        RECT -3.040 -24.705 -2.750 -24.660 ;
        RECT -0.940 -24.705 -0.650 -24.660 ;
        RECT 0.630 -24.705 0.920 -24.660 ;
        RECT 8.800 -24.750 12.100 -24.400 ;
        RECT -7.350 -25.100 -6.950 -25.050 ;
        RECT -8.950 -25.450 -6.950 -25.100 ;
        RECT -6.370 -25.110 -6.080 -25.010 ;
        RECT -2.645 -24.860 -2.355 -24.815 ;
        RECT -1.455 -24.860 -1.165 -24.815 ;
        RECT 1.065 -24.860 1.355 -24.815 ;
        RECT 10.400 -24.850 12.100 -24.750 ;
        RECT -2.645 -25.000 1.355 -24.860 ;
        RECT -2.645 -25.045 -2.355 -25.000 ;
        RECT -1.455 -25.045 -1.165 -25.000 ;
        RECT 1.065 -25.045 1.355 -25.000 ;
        RECT -6.370 -25.410 -4.490 -25.110 ;
        RECT -8.950 -30.350 -8.550 -25.450 ;
        RECT -7.350 -25.500 -6.950 -25.450 ;
        RECT -4.720 -25.700 -4.490 -25.410 ;
        RECT -2.260 -25.700 -1.980 -25.410 ;
        RECT 8.000 -25.450 8.750 -25.100 ;
        RECT 8.000 -25.550 8.300 -25.450 ;
        RECT -4.720 -26.000 -1.980 -25.700 ;
        RECT 6.250 -25.850 8.300 -25.550 ;
        RECT -8.950 -30.750 11.850 -30.350 ;
        RECT -5.220 -33.150 -4.930 -33.105 ;
        RECT -3.360 -33.150 -3.070 -33.105 ;
        RECT -0.580 -33.150 -0.290 -33.105 ;
        RECT -5.220 -33.290 -0.290 -33.150 ;
        RECT -5.220 -33.335 -4.930 -33.290 ;
        RECT -3.360 -33.335 -3.070 -33.290 ;
        RECT -0.580 -33.335 -0.290 -33.290 ;
        RECT 6.750 -33.330 9.050 -32.980 ;
        RECT -11.200 -34.100 -10.400 -33.700 ;
        RECT -6.750 -33.980 -3.600 -33.580 ;
        RECT -0.580 -33.830 -0.290 -33.785 ;
        RECT -2.825 -33.970 -0.290 -33.830 ;
        RECT -11.200 -50.100 -10.800 -34.100 ;
        RECT -8.050 -38.930 -7.600 -38.880 ;
        RECT -8.450 -39.280 -7.600 -38.930 ;
        RECT -8.050 -39.330 -7.600 -39.280 ;
        RECT -6.750 -40.830 -6.400 -33.980 ;
        RECT -2.825 -34.125 -2.610 -33.970 ;
        RECT -0.580 -34.015 -0.290 -33.970 ;
        RECT -4.760 -34.170 -4.470 -34.125 ;
        RECT -2.900 -34.170 -2.610 -34.125 ;
        RECT -1.980 -34.130 -1.690 -34.125 ;
        RECT -4.760 -34.310 -2.610 -34.170 ;
        RECT -4.760 -34.355 -4.470 -34.310 ;
        RECT -2.900 -34.355 -2.610 -34.310 ;
        RECT -2.050 -34.170 -1.550 -34.130 ;
        RECT 1.280 -34.170 1.570 -34.125 ;
        RECT -2.050 -34.310 1.570 -34.170 ;
        RECT -2.050 -34.580 -1.550 -34.310 ;
        RECT 1.280 -34.355 1.570 -34.310 ;
        RECT 4.700 -36.580 5.050 -33.730 ;
        RECT -2.650 -36.930 5.050 -36.580 ;
        RECT -2.650 -38.580 -2.300 -36.930 ;
        RECT -2.650 -38.930 0.250 -38.580 ;
        RECT -0.700 -39.780 -0.350 -39.430 ;
        RECT -0.100 -39.480 0.250 -38.930 ;
        RECT 4.550 -39.350 4.850 -38.680 ;
        RECT -0.200 -39.730 0.350 -39.480 ;
        RECT 4.550 -39.740 7.500 -39.350 ;
        RECT 4.850 -39.750 7.500 -39.740 ;
        RECT -9.400 -41.130 -6.400 -40.830 ;
        RECT -2.650 -40.130 -0.350 -39.780 ;
        RECT -9.400 -43.280 -9.050 -41.130 ;
        RECT -2.650 -41.830 -2.300 -40.130 ;
        RECT 8.700 -41.630 9.050 -33.330 ;
        RECT 11.450 -39.350 11.850 -30.750 ;
        RECT 10.650 -39.750 11.850 -39.350 ;
        RECT -6.400 -42.180 -2.300 -41.830 ;
        RECT 4.350 -41.980 9.050 -41.630 ;
        RECT -6.400 -43.230 -6.050 -42.180 ;
        RECT -9.400 -43.630 -7.350 -43.280 ;
        RECT -6.400 -43.630 -4.950 -43.230 ;
        RECT -3.410 -43.520 -3.120 -43.475 ;
        RECT -0.150 -43.520 0.350 -43.180 ;
        RECT -3.410 -43.660 0.350 -43.520 ;
        RECT -3.410 -43.705 -3.120 -43.660 ;
        RECT -0.150 -43.680 0.350 -43.660 ;
        RECT 0.770 -43.520 1.060 -43.475 ;
        RECT 2.630 -43.520 2.920 -43.475 ;
        RECT 0.770 -43.660 2.920 -43.520 ;
        RECT -0.150 -43.705 0.140 -43.680 ;
        RECT 0.770 -43.705 1.060 -43.660 ;
        RECT 2.630 -43.705 2.920 -43.660 ;
        RECT -1.550 -43.860 -1.260 -43.815 ;
        RECT 0.770 -43.860 0.985 -43.705 ;
        RECT -1.550 -44.000 0.985 -43.860 ;
        RECT -1.550 -44.045 -1.260 -44.000 ;
        RECT 1.750 -44.030 2.150 -43.830 ;
        RECT 4.350 -44.030 4.700 -41.980 ;
        RECT 19.250 -43.650 19.750 -12.500 ;
        RECT 30.150 -24.150 30.550 -8.100 ;
        RECT 31.900 -14.150 32.400 1.050 ;
        RECT 35.950 -0.700 36.350 1.050 ;
        RECT 39.300 -0.650 39.700 1.250 ;
        RECT 44.700 1.050 51.950 1.250 ;
        RECT 52.500 1.250 67.550 1.450 ;
        RECT 52.500 1.050 52.900 1.250 ;
        RECT 47.800 0.450 48.200 0.650 ;
        RECT 43.850 0.000 48.200 0.450 ;
        RECT 43.850 -0.650 44.300 0.000 ;
        RECT 47.800 -0.150 48.200 0.000 ;
        RECT 35.950 -1.150 38.000 -0.700 ;
        RECT 39.300 -1.150 41.600 -0.650 ;
        RECT 43.500 -1.150 44.450 -0.650 ;
        RECT 51.550 -0.700 51.950 1.050 ;
        RECT 54.900 -0.650 55.300 1.250 ;
        RECT 60.300 1.050 67.550 1.250 ;
        RECT 68.100 1.250 85.300 1.450 ;
        RECT 68.100 1.050 68.500 1.250 ;
        RECT 63.400 0.450 63.800 0.650 ;
        RECT 59.450 0.000 63.800 0.450 ;
        RECT 59.450 -0.650 59.900 0.000 ;
        RECT 63.400 -0.150 63.800 0.000 ;
        RECT 45.500 -1.150 48.900 -0.700 ;
        RECT 51.550 -1.150 53.600 -0.700 ;
        RECT 54.900 -1.150 57.200 -0.650 ;
        RECT 59.100 -1.150 60.050 -0.650 ;
        RECT 67.150 -0.700 67.550 1.050 ;
        RECT 70.500 -0.650 70.900 1.250 ;
        RECT 75.900 1.050 85.300 1.250 ;
        RECT 79.000 0.450 79.400 0.650 ;
        RECT 75.050 0.000 79.400 0.450 ;
        RECT 75.050 -0.650 75.500 0.000 ;
        RECT 79.000 -0.150 79.400 0.000 ;
        RECT 61.100 -1.150 64.500 -0.700 ;
        RECT 67.150 -1.150 69.200 -0.700 ;
        RECT 70.500 -1.150 72.800 -0.650 ;
        RECT 74.700 -1.150 75.650 -0.650 ;
        RECT 76.700 -1.150 80.100 -0.700 ;
        RECT 45.500 -2.250 45.900 -1.150 ;
        RECT 33.400 -2.650 45.900 -2.250 ;
        RECT 47.800 -2.250 48.200 -1.850 ;
        RECT 61.100 -2.250 61.500 -1.150 ;
        RECT 47.800 -2.650 61.500 -2.250 ;
        RECT 63.400 -2.250 63.800 -1.850 ;
        RECT 76.700 -2.250 77.100 -1.150 ;
        RECT 63.400 -2.650 77.100 -2.250 ;
        RECT 79.000 -2.250 79.400 -1.850 ;
        RECT 79.000 -2.650 83.800 -2.250 ;
        RECT 33.400 -10.450 33.900 -2.650 ;
        RECT 47.800 -3.050 48.200 -2.650 ;
        RECT 63.400 -3.050 63.800 -2.650 ;
        RECT 79.000 -3.050 79.400 -2.650 ;
        RECT 50.650 -10.450 51.050 -10.050 ;
        RECT 66.250 -10.450 66.650 -10.050 ;
        RECT 83.300 -10.450 83.800 -2.650 ;
        RECT 33.400 -10.850 51.050 -10.450 ;
        RECT 50.650 -11.250 51.050 -10.850 ;
        RECT 52.950 -10.850 66.650 -10.450 ;
        RECT 52.950 -11.950 53.350 -10.850 ;
        RECT 66.250 -11.250 66.650 -10.850 ;
        RECT 68.550 -10.850 83.800 -10.450 ;
        RECT 68.550 -11.950 68.950 -10.850 ;
        RECT 49.950 -12.400 53.350 -11.950 ;
        RECT 54.400 -12.450 55.350 -11.950 ;
        RECT 57.250 -12.450 59.550 -11.950 ;
        RECT 60.850 -12.400 62.900 -11.950 ;
        RECT 65.550 -12.400 68.950 -11.950 ;
        RECT 50.650 -13.100 51.050 -12.950 ;
        RECT 54.550 -13.100 55.000 -12.450 ;
        RECT 50.650 -13.550 55.000 -13.100 ;
        RECT 50.650 -13.750 51.050 -13.550 ;
        RECT 31.900 -14.350 54.150 -14.150 ;
        RECT 59.150 -14.350 59.550 -12.450 ;
        RECT 62.500 -14.150 62.900 -12.400 ;
        RECT 70.000 -12.450 70.950 -11.950 ;
        RECT 72.850 -12.450 75.150 -11.950 ;
        RECT 76.450 -12.400 78.500 -11.950 ;
        RECT 66.250 -13.100 66.650 -12.950 ;
        RECT 70.150 -13.100 70.600 -12.450 ;
        RECT 66.250 -13.550 70.600 -13.100 ;
        RECT 66.250 -13.750 66.650 -13.550 ;
        RECT 61.550 -14.350 61.950 -14.150 ;
        RECT 31.900 -14.550 61.950 -14.350 ;
        RECT 62.500 -14.350 69.750 -14.150 ;
        RECT 74.750 -14.350 75.150 -12.450 ;
        RECT 78.100 -14.150 78.500 -12.400 ;
        RECT 84.800 -14.150 85.300 1.050 ;
        RECT 77.150 -14.350 77.550 -14.150 ;
        RECT 62.500 -14.550 77.550 -14.350 ;
        RECT 78.100 -14.550 85.300 -14.150 ;
        RECT 47.100 -20.350 47.500 -14.550 ;
        RECT 53.750 -14.750 61.950 -14.550 ;
        RECT 53.750 -14.950 54.150 -14.750 ;
        RECT 61.550 -14.950 61.950 -14.750 ;
        RECT 69.350 -14.750 77.550 -14.550 ;
        RECT 69.350 -14.950 69.750 -14.750 ;
        RECT 77.150 -14.950 77.550 -14.750 ;
        RECT 52.950 -15.800 53.350 -15.300 ;
        RECT 56.050 -15.700 56.450 -15.200 ;
        RECT 59.150 -15.700 59.550 -15.200 ;
        RECT 63.850 -15.800 64.250 -15.300 ;
        RECT 68.550 -15.800 68.950 -15.300 ;
        RECT 71.650 -15.700 72.050 -15.200 ;
        RECT 74.750 -15.700 75.150 -15.200 ;
        RECT 79.450 -15.800 79.850 -15.300 ;
        RECT 86.300 -16.650 86.800 3.550 ;
        RECT 78.650 -17.050 86.800 -16.650 ;
        RECT 47.100 -20.750 58.450 -20.350 ;
        RECT 58.050 -21.800 58.450 -20.750 ;
        RECT 58.050 -21.810 60.150 -21.800 ;
        RECT 58.050 -22.170 60.480 -21.810 ;
        RECT 61.100 -21.850 61.350 -20.850 ;
        RECT 62.750 -21.850 67.350 -21.700 ;
        RECT 61.100 -22.050 67.350 -21.850 ;
        RECT 61.185 -22.060 67.350 -22.050 ;
        RECT 58.050 -22.200 60.150 -22.170 ;
        RECT 62.750 -22.200 67.350 -22.060 ;
        RECT 30.150 -24.550 32.600 -24.150 ;
        RECT 32.200 -35.750 32.600 -24.550 ;
        RECT 66.850 -25.650 67.350 -22.200 ;
        RECT 72.960 -25.120 73.250 -25.075 ;
        RECT 75.060 -25.120 75.350 -25.075 ;
        RECT 76.630 -25.120 76.920 -25.075 ;
        RECT 72.960 -25.260 76.920 -25.120 ;
        RECT 72.960 -25.305 73.250 -25.260 ;
        RECT 75.060 -25.305 75.350 -25.260 ;
        RECT 76.630 -25.305 76.920 -25.260 ;
        RECT 73.355 -25.460 73.645 -25.415 ;
        RECT 74.545 -25.460 74.835 -25.415 ;
        RECT 77.065 -25.460 77.355 -25.415 ;
        RECT 73.355 -25.600 77.355 -25.460 ;
        RECT 73.355 -25.645 73.645 -25.600 ;
        RECT 74.545 -25.645 74.835 -25.600 ;
        RECT 77.065 -25.645 77.355 -25.600 ;
        RECT 65.100 -25.950 68.300 -25.650 ;
        RECT 46.850 -26.500 47.250 -26.000 ;
        RECT 47.550 -26.150 47.950 -26.050 ;
        RECT 49.350 -26.150 49.750 -26.050 ;
        RECT 47.550 -26.700 49.750 -26.150 ;
        RECT 47.550 -26.850 47.950 -26.700 ;
        RECT 49.350 -26.850 49.750 -26.700 ;
        RECT 39.200 -29.750 39.600 -26.850 ;
        RECT 42.950 -27.750 45.150 -27.250 ;
        RECT 42.950 -27.850 43.350 -27.750 ;
        RECT 44.750 -27.850 45.150 -27.750 ;
        RECT 48.450 -27.850 50.650 -27.250 ;
        RECT 52.350 -29.750 52.750 -26.050 ;
        RECT 53.050 -29.750 53.450 -26.900 ;
        RECT 65.100 -27.650 65.400 -25.950 ;
        RECT 67.900 -26.050 68.300 -25.950 ;
        RECT 73.650 -26.200 74.150 -25.850 ;
        RECT 71.000 -26.550 74.150 -26.200 ;
        RECT 71.000 -26.750 71.550 -26.550 ;
        RECT 79.300 -26.650 87.500 -26.150 ;
        RECT 65.100 -27.950 69.050 -27.650 ;
        RECT 39.200 -30.150 53.450 -29.750 ;
        RECT 68.750 -30.000 69.050 -27.950 ;
        RECT 81.400 -28.950 81.900 -27.800 ;
        RECT 77.850 -29.200 81.900 -28.950 ;
        RECT 71.560 -29.320 71.850 -29.275 ;
        RECT 73.660 -29.320 73.950 -29.275 ;
        RECT 75.230 -29.320 75.520 -29.275 ;
        RECT 71.560 -29.460 75.520 -29.320 ;
        RECT 71.560 -29.505 71.850 -29.460 ;
        RECT 73.660 -29.505 73.950 -29.460 ;
        RECT 75.230 -29.505 75.520 -29.460 ;
        RECT 71.050 -30.000 71.450 -29.650 ;
        RECT 71.955 -29.660 72.245 -29.615 ;
        RECT 73.145 -29.660 73.435 -29.615 ;
        RECT 75.665 -29.660 75.955 -29.615 ;
        RECT 71.955 -29.800 75.955 -29.660 ;
        RECT 71.955 -29.845 72.245 -29.800 ;
        RECT 73.145 -29.845 73.435 -29.800 ;
        RECT 75.665 -29.845 75.955 -29.800 ;
        RECT 68.750 -30.300 71.450 -30.000 ;
        RECT 72.350 -30.550 72.750 -29.950 ;
        RECT 70.000 -30.800 72.750 -30.550 ;
        RECT 77.850 -30.000 78.300 -29.200 ;
        RECT 77.850 -30.750 78.350 -30.000 ;
        RECT 41.450 -32.500 46.850 -32.000 ;
        RECT 37.950 -33.550 38.350 -33.050 ;
        RECT 38.650 -33.250 39.050 -33.100 ;
        RECT 40.450 -33.250 40.850 -33.100 ;
        RECT 38.650 -33.750 40.850 -33.250 ;
        RECT 38.650 -33.900 39.050 -33.750 ;
        RECT 40.450 -33.900 40.850 -33.750 ;
        RECT 38.650 -36.450 39.050 -36.300 ;
        RECT 40.450 -36.450 40.850 -36.300 ;
        RECT 38.650 -36.950 40.850 -36.450 ;
        RECT 38.650 -37.100 39.050 -36.950 ;
        RECT 40.450 -37.100 40.850 -36.950 ;
        RECT 41.450 -37.500 41.950 -32.500 ;
        RECT 43.450 -33.450 43.850 -33.250 ;
        RECT 45.250 -33.450 45.650 -33.250 ;
        RECT 43.450 -33.950 45.650 -33.450 ;
        RECT 43.450 -34.100 43.850 -33.950 ;
        RECT 45.250 -34.100 45.650 -33.950 ;
        RECT 46.350 -35.650 46.850 -32.500 ;
        RECT 47.300 -33.750 47.700 -33.250 ;
        RECT 49.100 -33.750 49.500 -33.250 ;
        RECT 51.800 -33.700 52.200 -33.200 ;
        RECT 52.500 -33.300 52.900 -33.150 ;
        RECT 54.300 -33.300 54.700 -33.150 ;
        RECT 47.300 -34.250 49.500 -33.750 ;
        RECT 52.500 -33.800 54.700 -33.300 ;
        RECT 52.500 -33.950 52.900 -33.800 ;
        RECT 54.300 -33.950 54.700 -33.800 ;
        RECT 47.300 -34.400 47.700 -34.250 ;
        RECT 49.100 -34.400 49.500 -34.250 ;
        RECT 43.850 -36.150 45.250 -35.650 ;
        RECT 46.350 -36.150 49.100 -35.650 ;
        RECT 52.500 -36.500 52.900 -36.350 ;
        RECT 54.300 -36.500 54.700 -36.350 ;
        RECT 52.500 -37.000 54.700 -36.500 ;
        RECT 52.500 -37.150 52.900 -37.000 ;
        RECT 54.300 -37.150 54.700 -37.000 ;
        RECT 66.750 -37.350 67.250 -33.050 ;
        RECT 70.000 -34.050 70.500 -30.800 ;
        RECT 80.900 -30.900 81.400 -30.500 ;
        RECT 87.000 -34.050 87.500 -26.650 ;
        RECT 70.000 -34.550 87.500 -34.050 ;
        RECT 72.960 -36.820 73.250 -36.775 ;
        RECT 75.060 -36.820 75.350 -36.775 ;
        RECT 76.630 -36.820 76.920 -36.775 ;
        RECT 72.960 -36.960 76.920 -36.820 ;
        RECT 72.960 -37.005 73.250 -36.960 ;
        RECT 75.060 -37.005 75.350 -36.960 ;
        RECT 76.630 -37.005 76.920 -36.960 ;
        RECT 73.355 -37.160 73.645 -37.115 ;
        RECT 74.545 -37.160 74.835 -37.115 ;
        RECT 77.065 -37.160 77.355 -37.115 ;
        RECT 73.355 -37.300 77.355 -37.160 ;
        RECT 73.355 -37.345 73.645 -37.300 ;
        RECT 74.545 -37.345 74.835 -37.300 ;
        RECT 77.065 -37.345 77.355 -37.300 ;
        RECT 39.050 -38.000 41.950 -37.500 ;
        RECT 52.900 -38.050 54.700 -37.550 ;
        RECT 32.600 -39.450 33.450 -39.100 ;
        RECT 39.350 -39.250 40.150 -38.550 ;
        RECT 32.600 -41.100 33.100 -39.450 ;
        RECT 39.550 -42.450 39.950 -39.250 ;
        RECT 54.300 -40.000 54.700 -38.050 ;
        RECT 65.100 -37.650 68.300 -37.350 ;
        RECT 65.100 -39.350 65.400 -37.650 ;
        RECT 67.900 -37.750 68.300 -37.650 ;
        RECT 73.650 -37.900 74.150 -37.550 ;
        RECT 71.000 -38.250 74.150 -37.900 ;
        RECT 71.000 -38.450 71.550 -38.250 ;
        RECT 79.300 -38.350 87.500 -37.850 ;
        RECT 65.100 -39.650 69.050 -39.350 ;
        RECT 68.750 -41.700 69.050 -39.650 ;
        RECT 81.400 -39.850 82.450 -39.350 ;
        RECT 81.400 -40.650 81.900 -39.850 ;
        RECT 77.850 -40.900 81.900 -40.650 ;
        RECT 71.560 -41.020 71.850 -40.975 ;
        RECT 73.660 -41.020 73.950 -40.975 ;
        RECT 75.230 -41.020 75.520 -40.975 ;
        RECT 71.560 -41.160 75.520 -41.020 ;
        RECT 71.560 -41.205 71.850 -41.160 ;
        RECT 73.660 -41.205 73.950 -41.160 ;
        RECT 75.230 -41.205 75.520 -41.160 ;
        RECT 71.050 -41.700 71.450 -41.350 ;
        RECT 71.955 -41.360 72.245 -41.315 ;
        RECT 73.145 -41.360 73.435 -41.315 ;
        RECT 75.665 -41.360 75.955 -41.315 ;
        RECT 71.955 -41.500 75.955 -41.360 ;
        RECT 71.955 -41.545 72.245 -41.500 ;
        RECT 73.145 -41.545 73.435 -41.500 ;
        RECT 75.665 -41.545 75.955 -41.500 ;
        RECT 68.750 -42.000 71.450 -41.700 ;
        RECT 72.350 -42.250 72.750 -41.650 ;
        RECT 39.550 -42.520 41.000 -42.450 ;
        RECT 70.000 -42.500 72.750 -42.250 ;
        RECT 77.850 -41.700 78.300 -40.900 ;
        RECT 77.850 -42.450 78.350 -41.700 ;
        RECT 39.550 -42.770 42.965 -42.520 ;
        RECT 39.550 -42.850 41.000 -42.770 ;
        RECT 1.750 -44.330 4.700 -44.030 ;
        RECT 5.050 -44.080 6.700 -43.730 ;
        RECT 1.750 -44.380 2.950 -44.330 ;
        RECT 3.550 -44.380 4.700 -44.330 ;
        RECT -1.550 -44.540 -1.260 -44.495 ;
        RECT 1.230 -44.540 1.520 -44.495 ;
        RECT 3.090 -44.540 3.380 -44.495 ;
        RECT -1.550 -44.680 3.380 -44.540 ;
        RECT -1.550 -44.725 -1.260 -44.680 ;
        RECT 1.230 -44.725 1.520 -44.680 ;
        RECT 3.090 -44.725 3.380 -44.680 ;
        RECT 6.350 -44.880 6.700 -44.080 ;
        RECT 18.750 -44.150 19.750 -43.650 ;
        RECT 70.000 -45.750 70.500 -42.500 ;
        RECT 80.900 -42.600 81.400 -42.200 ;
        RECT 87.000 -45.750 87.500 -38.350 ;
        RECT 70.000 -46.250 87.500 -45.750 ;
        RECT 85.350 -50.100 85.850 -49.700 ;
        RECT -11.200 -50.500 85.850 -50.100 ;
      LAYER met2 ;
        RECT -2.050 -3.030 -1.550 -2.480 ;
        RECT -2.050 -4.180 -1.700 -3.030 ;
        RECT -5.200 -4.530 -1.700 -4.180 ;
        RECT -8.050 -7.280 -7.600 -7.230 ;
        RECT -5.200 -7.280 -4.850 -4.530 ;
        RECT -8.050 -7.630 -4.850 -7.280 ;
        RECT -8.050 -7.680 -7.600 -7.630 ;
        RECT -5.200 -9.580 -4.850 -7.630 ;
        RECT -5.200 -9.930 0.200 -9.580 ;
        RECT -0.150 -11.530 0.200 -9.930 ;
        RECT -0.150 -12.030 0.350 -11.530 ;
        RECT 81.400 -28.300 86.050 -27.800 ;
        RECT 85.550 -33.050 86.050 -28.300 ;
        RECT 66.750 -33.550 86.050 -33.050 ;
        RECT -2.050 -34.680 -1.550 -34.130 ;
        RECT -2.050 -35.830 -1.700 -34.680 ;
        RECT -5.200 -36.180 -1.700 -35.830 ;
        RECT -8.050 -38.930 -7.600 -38.880 ;
        RECT -5.200 -38.930 -4.850 -36.180 ;
        RECT -8.050 -39.280 -4.850 -38.930 ;
        RECT -8.050 -39.330 -7.600 -39.280 ;
        RECT -5.200 -41.230 -4.850 -39.280 ;
        RECT -5.200 -41.580 0.200 -41.230 ;
        RECT -0.150 -43.180 0.200 -41.580 ;
        RECT -0.150 -43.680 0.350 -43.180 ;
  END
END vco_adc2
END LIBRARY

