magic
tech sky130A
magscale 1 2
timestamp 1730530608
<< nwell >>
rect -410 310 20 640
rect 520 300 940 630
rect -610 -530 -440 -210
rect 180 -540 650 -210
rect 2640 -260 2940 -210
rect 2630 -270 2940 -260
rect 2640 -540 2940 -270
<< pwell >>
rect -410 60 60 260
rect 480 60 970 210
rect -610 -840 -390 -590
rect 120 -780 690 -630
rect 2610 -780 2940 -590
<< psubdiff >>
rect -350 170 -270 200
rect -350 130 -330 170
rect -290 130 -270 170
rect -350 100 -270 130
rect 2660 -660 2760 -640
rect -550 -710 -470 -680
rect -550 -750 -530 -710
rect -490 -750 -470 -710
rect 2660 -700 2690 -660
rect 2730 -700 2760 -660
rect 2660 -720 2760 -700
rect -550 -780 -470 -750
<< nsubdiff >>
rect -350 500 -270 530
rect -350 460 -330 500
rect -290 460 -270 500
rect -350 430 -270 460
rect -550 -350 -470 -320
rect -550 -390 -530 -350
rect -490 -390 -470 -350
rect -550 -420 -470 -390
rect 2680 -430 2780 -410
rect 2680 -470 2710 -430
rect 2750 -470 2780 -430
rect 2680 -490 2780 -470
<< psubdiffcont >>
rect -330 130 -290 170
rect -530 -750 -490 -710
rect 2690 -700 2730 -660
<< nsubdiffcont >>
rect -330 460 -290 500
rect -530 -390 -490 -350
rect 2710 -470 2750 -430
<< locali >>
rect 2420 570 2690 640
rect -350 500 -270 530
rect -350 460 -330 500
rect -290 460 -270 500
rect -350 430 -270 460
rect 470 290 980 370
rect -1590 170 -270 200
rect -1590 130 -1560 170
rect -1520 130 -330 170
rect -290 130 -270 170
rect -1590 100 -270 130
rect 680 170 790 200
rect 680 130 720 170
rect 760 130 790 170
rect 680 110 790 130
rect 715 -65 765 110
rect 560 -115 765 -65
rect 150 -220 480 -200
rect 150 -260 410 -220
rect 450 -260 480 -220
rect 150 -290 480 -260
rect -550 -350 -470 -320
rect -550 -390 -530 -350
rect -490 -390 -470 -350
rect 560 -370 610 -115
rect 2610 -120 2690 570
rect 2610 -160 2630 -120
rect 2670 -160 2690 -120
rect 2610 -180 2690 -160
rect -550 -420 -470 -390
rect 150 -420 610 -370
rect 150 -530 205 -420
rect 2680 -430 2780 -410
rect 2680 -470 2710 -430
rect 2750 -470 2780 -430
rect 2680 -490 2780 -470
rect -700 -570 -370 -530
rect -700 -1000 -640 -570
rect 0 -580 205 -530
rect 2490 -530 2500 -520
rect 2490 -570 2900 -530
rect 2490 -580 2500 -570
rect 2630 -600 2900 -570
rect 2660 -660 2760 -640
rect -550 -710 -470 -680
rect -550 -750 -530 -710
rect -490 -750 -470 -710
rect 2660 -700 2690 -660
rect 2730 -700 2760 -660
rect 2660 -720 2760 -700
rect -550 -780 -470 -750
rect 150 -840 680 -740
rect 2820 -1000 2900 -600
rect -700 -1080 2900 -1000
<< viali >>
rect -330 460 -290 500
rect 70 270 110 310
rect 1240 210 1280 250
rect -1560 130 -1520 170
rect -330 130 -290 170
rect 720 130 760 170
rect 2350 150 2390 190
rect 410 -260 450 -220
rect -530 -390 -490 -350
rect 2630 -160 2670 -120
rect 2070 -390 2110 -350
rect 2070 -470 2110 -430
rect 2710 -470 2750 -430
rect 710 -580 750 -540
rect 960 -610 1000 -570
rect 2070 -680 2110 -640
rect -530 -750 -490 -710
rect 2690 -700 2730 -660
<< metal1 >>
rect 490 540 980 640
rect -1160 500 -270 530
rect -1160 460 -330 500
rect -290 460 -270 500
rect -1160 430 -270 460
rect -1590 170 -1490 200
rect -1590 130 -1560 170
rect -1520 130 -1490 170
rect -1590 -680 -1490 130
rect -1160 -320 -1060 430
rect -500 310 140 330
rect -500 270 70 310
rect 110 270 140 310
rect -500 -70 -440 270
rect 60 250 140 270
rect 1210 250 1310 290
rect 1210 220 1240 250
rect 680 210 1240 220
rect 1280 210 1310 250
rect -350 170 -270 200
rect -350 130 -330 170
rect -290 130 -270 170
rect -350 100 -270 130
rect 680 170 1310 210
rect 680 130 720 170
rect 760 150 1310 170
rect 2340 190 3980 230
rect 2340 150 2350 190
rect 2390 150 3980 190
rect 760 130 790 150
rect 2340 130 3980 150
rect 680 110 790 130
rect 490 0 960 70
rect 2430 0 3380 80
rect -500 -130 290 -70
rect -550 -290 -380 -200
rect -550 -320 -470 -290
rect -1160 -350 -470 -320
rect -1160 -390 -530 -350
rect -490 -390 -470 -350
rect -1160 -420 -470 -390
rect 230 -540 290 -130
rect 2610 -120 2690 -100
rect 2610 -160 2630 -120
rect 2670 -160 2690 -120
rect 380 -220 690 -200
rect 380 -260 410 -220
rect 450 -260 690 -220
rect 380 -290 690 -260
rect 2610 -300 2690 -160
rect 2760 -330 2860 -130
rect 2050 -350 2860 -330
rect 2050 -390 2070 -350
rect 2110 -380 2860 -350
rect 2110 -390 2140 -380
rect 2050 -430 2140 -390
rect 2050 -470 2070 -430
rect 2110 -470 2140 -430
rect 690 -540 770 -470
rect 230 -580 710 -540
rect 750 -580 770 -540
rect 230 -600 770 -580
rect 950 -570 1030 -530
rect 950 -610 960 -570
rect 1000 -610 1030 -570
rect 950 -650 1030 -610
rect -1590 -710 -470 -680
rect -1590 -750 -530 -710
rect -490 -750 -470 -710
rect 480 -700 1030 -650
rect 2050 -540 2140 -470
rect 2680 -430 2780 -410
rect 2680 -470 2710 -430
rect 2750 -470 2780 -430
rect 2680 -490 2780 -470
rect 2050 -640 2150 -540
rect 2050 -680 2070 -640
rect 2110 -680 2150 -640
rect 2050 -690 2150 -680
rect 2660 -660 2760 -640
rect 2660 -700 2690 -660
rect 2730 -700 2760 -660
rect -1590 -780 -390 -750
rect -550 -840 -390 -780
rect 480 -1350 580 -700
rect 2660 -720 2760 -700
rect 3290 -750 3380 0
rect 2610 -840 3380 -750
rect 3880 -1350 3980 130
rect 480 -1450 3980 -1350
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -402 0 1 -792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_2  sky130_fd_sc_hd__dfxbp_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 678 0 1 -792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 958 0 1 48
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 38 0 1 48
box -38 -48 498 592
<< labels >>
rlabel metal1 230 -70 230 -70 1 clk
port 1 n
rlabel locali 180 -580 180 -580 5 Q_N_buf
rlabel locali -660 -530 -660 -530 1 Q_N
rlabel metal1 2580 230 2580 230 1 D
rlabel locali 680 290 680 290 5 clkinv
rlabel metal1 2810 -130 2810 -130 1 clkDiv2
port 2 n
rlabel metal1 -1540 200 -1540 200 1 GND
port 4 n
rlabel metal1 -1100 530 -1100 530 1 VDDA
port 3 n
<< end >>
