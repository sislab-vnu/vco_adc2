magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect 730 650 5670 730
rect 690 390 5670 650
rect 920 -120 4190 -70
rect 690 -410 4190 -120
<< pwell >>
rect 3114 162 3228 314
rect 1104 -616 1236 -464
<< psubdiff >>
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 3140 188 3202 224
rect 1130 -523 1210 -490
rect 1130 -557 1153 -523
rect 1187 -557 1210 -523
rect 1130 -590 1210 -557
<< nsubdiff >>
rect 3150 567 3230 600
rect 3150 533 3173 567
rect 3207 533 3230 567
rect 3150 500 3230 533
rect 1180 -233 1260 -200
rect 1180 -267 1203 -233
rect 1237 -267 1260 -233
rect 1180 -300 1260 -267
<< psubdiffcont >>
rect 3156 224 3190 258
rect 1153 -557 1187 -523
<< nsubdiffcont >>
rect 3173 533 3207 567
rect 1203 -267 1237 -233
<< locali >>
rect 730 680 810 730
rect 3150 567 3230 600
rect 3150 533 3173 567
rect 3207 533 3230 567
rect 3150 500 3230 533
rect 1420 350 1650 460
rect 2260 350 2450 460
rect 3080 350 3290 460
rect 3960 350 4150 460
rect 4770 350 4920 460
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 5590 250 5890 320
rect 3140 188 3202 224
rect 5820 50 5890 250
rect 3700 -20 5890 50
rect 1020 -110 1570 -70
rect 1180 -233 1260 -110
rect 1180 -267 1203 -233
rect 1237 -267 1260 -233
rect 1180 -300 1260 -267
rect 3700 -400 3770 -20
rect 3990 -253 4030 -250
rect 3990 -287 3993 -253
rect 4027 -287 4030 -253
rect 3990 -290 4030 -287
rect 760 -413 800 -410
rect 760 -447 763 -413
rect 797 -447 800 -413
rect 760 -450 800 -447
rect 2930 -450 3420 -400
rect 3590 -450 3770 -400
rect 3900 -403 3940 -400
rect 3900 -437 3903 -403
rect 3937 -437 3940 -403
rect 3900 -440 3940 -437
rect 1130 -523 1210 -490
rect 3520 -493 3560 -490
rect 1130 -557 1153 -523
rect 1187 -557 1210 -523
rect 3520 -527 3523 -493
rect 3557 -527 3560 -493
rect 3520 -530 3560 -527
rect 1130 -590 1210 -557
<< viali >>
rect 3173 533 3207 567
rect 810 368 844 402
rect 3156 224 3190 258
rect 948 -286 982 -252
rect 1203 -267 1237 -233
rect 3993 -287 4027 -253
rect 763 -447 797 -413
rect 1516 -444 1550 -410
rect 3903 -437 3937 -403
rect 1768 -500 1802 -466
rect 1153 -557 1187 -523
rect 3523 -527 3557 -493
<< metal1 >>
rect 190 630 750 730
rect 1460 630 1560 730
rect 2280 630 2380 730
rect 3100 630 3250 730
rect 3980 630 4070 730
rect 4800 630 4890 730
rect 190 -70 290 630
rect 3150 567 3230 630
rect 3150 533 3173 567
rect 3207 533 3230 567
rect 3150 500 3230 533
rect 746 440 886 464
rect 440 402 886 440
rect 440 370 810 402
rect 440 40 510 370
rect 746 368 810 370
rect 844 368 886 402
rect 746 350 886 368
rect 3140 258 3202 288
rect 3140 224 3156 258
rect 3190 224 3202 258
rect 3140 190 3202 224
rect 1460 90 1550 190
rect 2280 90 2370 190
rect 3100 90 3250 190
rect 3980 90 4070 190
rect 440 -30 1410 40
rect 190 -170 750 -70
rect 934 -252 994 -202
rect 934 -286 948 -252
rect 982 -286 994 -252
rect 934 -372 994 -286
rect 1180 -233 1260 -200
rect 1180 -267 1203 -233
rect 1237 -267 1260 -233
rect 1180 -300 1260 -267
rect 740 -390 820 -380
rect 440 -413 820 -390
rect 440 -447 763 -413
rect 797 -447 820 -413
rect 440 -460 820 -447
rect 936 -392 994 -372
rect 1340 -330 1410 -30
rect 2960 -170 3340 -70
rect 3610 -170 3870 -70
rect 3970 -250 4050 -220
rect 3970 -253 4370 -250
rect 3970 -287 3993 -253
rect 4027 -287 4370 -253
rect 3970 -320 4370 -287
rect 1340 -338 1570 -330
rect 936 -452 1312 -392
rect 1340 -400 1572 -338
rect 740 -470 820 -460
rect 1130 -523 1210 -490
rect 1130 -557 1153 -523
rect 1187 -557 1210 -523
rect 1130 -610 1210 -557
rect 1266 -510 1312 -452
rect 1502 -410 1572 -400
rect 1502 -444 1516 -410
rect 1550 -444 1572 -410
rect 1502 -468 1572 -444
rect 3810 -403 3960 -390
rect 3810 -437 3903 -403
rect 3937 -437 3960 -403
rect 1758 -466 1814 -452
rect 1758 -500 1768 -466
rect 1802 -500 1814 -466
rect 3810 -460 3960 -437
rect 3810 -480 3870 -460
rect 1758 -510 1814 -500
rect 1266 -570 1814 -510
rect 3460 -493 3870 -480
rect 3460 -527 3523 -493
rect 3557 -527 3870 -493
rect 3460 -540 3870 -527
rect 4692 -610 4787 147
rect 4800 90 4890 190
rect 1090 -710 1490 -610
rect 2960 -710 3340 -610
rect 3610 -710 3870 -610
rect 4130 -615 4787 -610
rect 4093 -710 4787 -615
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0
timestamp 1729593089
transform 1 0 728 0 1 -662
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1729593089
transform 1 0 1488 0 1 -662
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_0
timestamp 1729593089
transform 1 0 728 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_1
timestamp 1729593089
transform 1 0 1548 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_2
timestamp 1729593089
transform 1 0 2368 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_3
timestamp 1729593089
transform 1 0 3248 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_4
timestamp 1729593089
transform 1 0 4068 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  sky130_fd_sc_hd__dlygate4sd3_1_5
timestamp 1729593089
transform 1 0 4888 0 1 138
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1729593089
transform 1 0 3868 0 1 -662
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1729593089
transform 1 0 3338 0 1 -662
box -38 -48 314 592
<< labels >>
rlabel locali s 5770 320 5770 320 4 CLK_dly
rlabel metal1 s 3640 -480 3640 -480 4 FBack_inv
rlabel locali s 1530 460 1530 460 4 DL1
rlabel locali s 2370 460 2370 460 4 DL2
rlabel locali s 3250 460 3250 460 4 DL3
rlabel locali s 4060 460 4060 460 4 DL4
rlabel locali s 4870 460 4870 460 4 DL5
rlabel metal1 s 490 440 490 440 4 CLK
rlabel locali s 3140 -400 3140 -400 4 Dout
rlabel metal1 s 4230 -250 4230 -250 4 FBack
rlabel metal1 s 540 -390 540 -390 4 D
rlabel metal1 s 4470 -610 4470 -610 4 GND
rlabel metal1 s 620 730 620 730 4 VCCD
<< end >>
