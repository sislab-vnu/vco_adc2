magic
tech sky130A
timestamp 1726649572
<< locali >>
rect 110 670 590 710
rect 110 400 150 670
rect 480 420 520 670
rect 550 430 590 670
rect 200 -105 240 200
rect 270 -105 310 200
rect 640 -105 680 70
rect 200 -145 680 -105
use n_lk  n_lk_0
timestamp 1726647885
transform -1 0 200 0 -1 400
box -130 -40 200 280
use p_lk  p_lk_0
timestamp 1726647848
transform 1 0 590 0 1 40
box -130 -40 200 490
<< labels >>
rlabel locali 365 710 365 710 1 add_pwr
rlabel locali 385 -105 385 -105 1 input_R
<< end >>
