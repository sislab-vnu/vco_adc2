magic
tech sky130A
magscale 1 2
timestamp 1729753075
<< locali >>
rect 1350 3520 3140 3660
rect 1350 0 1550 3520
rect 1350 -100 1400 0
rect 1500 -100 1550 0
rect -4740 -1610 -4370 -1600
rect -4740 -1794 -4646 -1610
rect -4462 -1630 -4370 -1610
rect 1350 -1630 1550 -100
rect -4462 -1794 1550 -1630
rect -4740 -1830 1550 -1794
rect -4740 -3890 -4370 -1830
rect -3300 -2860 -3200 -2830
rect -3300 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3300 -2920 -3200 -2900
rect 1350 -3230 1550 -1830
rect 19560 -2490 21710 -2480
rect 19560 -2530 19580 -2490
rect 19620 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 19560 -2550 21710 -2530
rect 18400 -3082 18470 -2660
rect 1350 -3370 5590 -3230
rect 1350 -3410 5520 -3370
rect 5560 -3410 5590 -3370
rect 1350 -3430 5590 -3410
rect -4740 -3930 -4460 -3890
rect -4420 -3930 -4370 -3890
rect -4740 -3950 -4370 -3930
rect 390 -4850 570 -4820
rect 390 -4890 500 -4850
rect 540 -4890 570 -4850
rect 390 -4920 570 -4890
rect 14710 -7240 14900 -7200
rect 14710 -7270 15490 -7240
rect 14710 -7320 14780 -7270
rect 14830 -7320 15490 -7270
rect 14710 -7380 14900 -7320
rect 19080 -9260 19180 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 19180 -9260
rect 19080 -9330 19180 -9300
<< viali >>
rect 540 7650 580 7690
rect 1630 7650 1670 7690
rect 2720 7650 2760 7690
rect 4640 7650 4680 7690
rect 6540 7650 6580 7690
rect 7630 7650 7670 7690
rect 8720 7650 8760 7690
rect 10640 7650 10680 7690
rect 12540 7650 12580 7690
rect 13630 7650 13670 7690
rect 14720 7650 14760 7690
rect 17970 7640 18030 7700
rect 6400 1000 6440 1040
rect 7490 1000 7530 1040
rect 8580 1000 8620 1040
rect 10480 1000 10520 1040
rect 12400 1000 12440 1040
rect 13490 1000 13530 1040
rect 14580 1000 14620 1040
rect 16480 1000 16520 1040
rect 17980 990 18040 1050
rect 1400 -100 1500 0
rect -4646 -1794 -4462 -1610
rect -3270 -2900 -3230 -2860
rect 19580 -2530 19620 -2490
rect 21650 -2530 21690 -2490
rect 18354 -3266 18538 -3082
rect 5520 -3410 5560 -3370
rect -4460 -3930 -4420 -3890
rect 500 -4890 540 -4850
rect 5460 -6320 5560 -6220
rect 14780 -7320 14830 -7270
rect 19110 -9300 19150 -9260
rect 19370 -9640 19470 -9540
<< metal1 >>
rect -1380 8050 -1180 8110
rect -1380 7950 -1340 8050
rect -1240 7950 -1180 8050
rect 11760 7980 11770 8080
rect 11870 7980 11880 8080
rect -1380 7910 -1180 7950
rect -1340 4930 -1330 5030
rect -1230 4930 -1220 5030
rect 14670 4880 14680 4980
rect 14780 4880 14790 4980
rect 1968 4462 1978 4646
rect 2162 4462 2172 4646
rect 3730 4050 3750 4150
rect 3840 4070 3850 4130
rect 3910 4070 3920 4130
rect -3390 1560 -1760 1660
rect -4658 -1610 -4450 -1604
rect -4658 -1794 -4646 -1610
rect -4462 -1794 -4450 -1610
rect -4658 -1800 -4450 -1794
rect -3390 -2830 -3300 1560
rect 13640 680 13740 710
rect 1350 0 15230 50
rect 1350 -100 1400 0
rect 1500 -100 15230 0
rect 1350 -150 15230 -100
rect 6380 -720 6460 -690
rect 13640 -1070 13740 -690
rect -3390 -2860 -3200 -2830
rect -3390 -2900 -3270 -2860
rect -3230 -2900 -3200 -2860
rect -3390 -2920 -3200 -2900
rect -3650 -3056 -3450 -3010
rect -3650 -3060 -3060 -3056
rect -3650 -3160 -3600 -3060
rect -3500 -3156 -3060 -3060
rect -3500 -3160 -3450 -3156
rect -3650 -3210 -3450 -3160
rect 5500 -3370 5570 -3350
rect 5500 -3410 5520 -3370
rect 5560 -3410 5570 -3370
rect 5500 -3430 5570 -3410
rect -3350 -3600 -3150 -3550
rect -3350 -3700 -3300 -3600
rect -3200 -3700 -3150 -3600
rect -3350 -3750 -3150 -3700
rect -4470 -3890 -3160 -3870
rect -4470 -3930 -4460 -3890
rect -4420 -3930 -3160 -3890
rect -4470 -3950 -3160 -3930
rect -70 -3970 60 -3960
rect -70 -4030 -10 -3970
rect 50 -4030 60 -3970
rect -70 -4040 60 -4030
rect 470 -4850 570 -4820
rect 470 -4890 500 -4850
rect 540 -4890 570 -4850
rect 470 -12490 570 -4890
rect 5200 -5980 5210 -5930
rect 5160 -6030 5210 -5980
rect 5310 -5980 5320 -5930
rect 5310 -6030 5440 -5980
rect 5160 -6080 5440 -6030
rect 6580 -6210 6680 -6190
rect 5448 -6220 5572 -6214
rect 5448 -6320 5460 -6220
rect 5560 -6320 5572 -6220
rect 6568 -6302 6578 -6210
rect 6670 -6302 6680 -6210
rect 5448 -6326 5572 -6320
rect 6580 -6420 6680 -6302
rect 14710 -7260 14900 -7200
rect 14710 -7330 14770 -7260
rect 14840 -7330 14900 -7260
rect 14710 -7380 14900 -7330
rect 15030 -8286 15230 -150
rect 20740 -1450 20750 -1350
rect 20850 -1450 20860 -1350
rect 20740 -1520 20860 -1450
rect 15676 -1886 15686 -1794
rect 15778 -1886 15788 -1794
rect 19560 -2490 19640 -2470
rect 19560 -2530 19580 -2490
rect 19620 -2530 19640 -2490
rect 19560 -2550 19640 -2530
rect 21610 -2490 21710 -2480
rect 21610 -2530 21650 -2490
rect 21690 -2530 21710 -2490
rect 15480 -2640 15800 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2690 15800 -2640
rect 15560 -2700 15580 -2690
rect 15480 -2720 15580 -2700
rect 19950 -2790 20150 -2740
rect 19950 -2890 20000 -2790
rect 20100 -2890 20150 -2790
rect 19950 -2940 20150 -2890
rect 18342 -3082 18550 -3076
rect 18342 -3266 18354 -3082
rect 18538 -3266 18550 -3082
rect 18342 -3272 18550 -3266
rect 15030 -8356 15570 -8286
rect 15030 -8370 15230 -8356
rect 18700 -8376 18800 -8360
rect 18540 -8380 18800 -8376
rect 18540 -8440 18720 -8380
rect 18780 -8440 18800 -8380
rect 18540 -8446 18800 -8440
rect 18700 -8460 18800 -8446
rect 19010 -9100 19150 -9000
rect 19250 -9100 19260 -9000
rect 21610 -9230 21710 -2530
rect 19080 -9260 21710 -9230
rect 19080 -9300 19110 -9260
rect 19150 -9300 21710 -9260
rect 19080 -9330 21710 -9300
rect 19358 -9540 19482 -9534
rect 19358 -9640 19370 -9540
rect 19470 -9640 19482 -9540
rect 19358 -9646 19482 -9640
rect 3630 -9900 3830 -9850
rect 3630 -10000 3680 -9900
rect 3780 -10000 3830 -9900
rect 3630 -10050 3830 -10000
rect 21610 -12490 21710 -9330
rect 470 -12590 21710 -12490
<< via1 >>
rect -1340 7950 -1240 8050
rect 11770 7980 11870 8080
rect -1330 4930 -1230 5030
rect 14680 4880 14780 4980
rect 1978 4462 2162 4646
rect 3850 4070 3910 4130
rect -4646 -1794 -4462 -1610
rect -3600 -3160 -3500 -3060
rect -3300 -3700 -3200 -3600
rect -10 -4030 50 -3970
rect 5210 -6030 5310 -5930
rect 5460 -6320 5560 -6220
rect 6578 -6302 6670 -6210
rect 14770 -7270 14840 -7260
rect 14770 -7320 14780 -7270
rect 14780 -7320 14830 -7270
rect 14830 -7320 14840 -7270
rect 14770 -7330 14840 -7320
rect 3870 -8260 3930 -8200
rect 20750 -1450 20850 -1350
rect 15686 -1886 15778 -1794
rect 15500 -2700 15560 -2640
rect 20000 -2890 20100 -2790
rect 18354 -3266 18538 -3082
rect 18720 -8440 18780 -8380
rect 19150 -9100 19250 -9000
rect 13720 -9310 13780 -9250
rect 19370 -9640 19470 -9540
rect 3680 -10000 3780 -9900
<< metal2 >>
rect -4738 -1610 -4370 8326
rect -3450 4738 -3082 8326
rect 11770 8080 11870 8090
rect -1340 8050 -1240 8060
rect 11770 7970 11870 7980
rect -1340 7940 -1240 7950
rect -1330 5030 -1230 5040
rect -1330 4920 -1230 4930
rect 14680 4980 14780 4990
rect 14680 4870 14780 4880
rect -3450 4646 2254 4738
rect -3450 4462 1978 4646
rect 2162 4462 2254 4646
rect -3450 4370 2254 4462
rect 3730 4140 3930 4150
rect 3730 4070 3750 4140
rect 3820 4130 3930 4140
rect 3820 4070 3850 4130
rect 3910 4070 3930 4130
rect 3730 4050 3930 4070
rect 20838 -230 21206 8326
rect -4738 -1794 -4646 -1610
rect -4462 -1794 -4370 -1610
rect -4738 -1886 -4370 -1794
rect 15594 -598 21206 -230
rect 15594 -1794 15870 -598
rect 20750 -1350 20850 -1340
rect 20750 -1460 20850 -1450
rect 15594 -1886 15686 -1794
rect 15778 -1886 15870 -1794
rect 15594 -1978 15870 -1886
rect 15480 -2640 15580 -2620
rect 15480 -2700 15500 -2640
rect 15560 -2700 15580 -2640
rect -3600 -3060 -3500 -3050
rect -3600 -3170 -3500 -3160
rect -3300 -3600 -3200 -3590
rect -3300 -3710 -3200 -3700
rect -20 -3970 1000 -3960
rect -20 -4030 -10 -3970
rect 50 -4030 1000 -3970
rect -20 -4040 1000 -4030
rect 920 -7670 1000 -4040
rect 4554 -5930 5360 -5880
rect 4554 -6030 5210 -5930
rect 5310 -6030 5360 -5930
rect 4554 -6080 5360 -6030
rect 4110 -6820 4210 -6810
rect 4110 -6930 4210 -6920
rect 920 -7750 3940 -7670
rect 3860 -8180 3940 -7750
rect 3850 -8200 3950 -8180
rect 3850 -8260 3870 -8200
rect 3930 -8260 3950 -8200
rect 3850 -8270 3950 -8260
rect 3680 -9900 3780 -9890
rect 3680 -10010 3780 -10000
rect 4554 -13570 4830 -6080
rect 6486 -6210 6762 -6118
rect 5460 -6220 5560 -6210
rect 5460 -6330 5560 -6320
rect 6486 -6302 6578 -6210
rect 6670 -6302 6762 -6210
rect 6486 -13570 6762 -6302
rect 15480 -6300 15580 -2700
rect 20000 -2790 20100 -2780
rect 20000 -2900 20100 -2890
rect 22402 -2990 22770 8326
rect 18262 -3082 22770 -2990
rect 18262 -3266 18354 -3082
rect 18538 -3266 22770 -3082
rect 18262 -3358 22770 -3266
rect 15480 -6400 19700 -6300
rect 14710 -7260 14900 -7200
rect 14710 -7330 14770 -7260
rect 14840 -7330 14900 -7260
rect 14710 -7379 14900 -7330
rect 9150 -8610 9250 -8600
rect 9150 -8720 9250 -8710
rect 13700 -9240 13800 -9220
rect 14750 -9240 14853 -7379
rect 19600 -8360 19700 -6400
rect 18700 -8380 19700 -8360
rect 18700 -8440 18720 -8380
rect 18780 -8440 19700 -8380
rect 18700 -8460 19700 -8440
rect 19150 -9000 19250 -8990
rect 19150 -9110 19250 -9100
rect 13700 -9250 14853 -9240
rect 13700 -9310 13720 -9250
rect 13780 -9310 14853 -9250
rect 13700 -9340 14853 -9310
rect 19370 -9540 19470 -9530
rect 19370 -9650 19470 -9640
<< via2 >>
rect -1340 7950 -1240 8050
rect 11770 7980 11870 8080
rect -1330 4930 -1230 5030
rect 14680 4880 14780 4980
rect 3750 4070 3820 4140
rect 20750 -1450 20850 -1350
rect -3600 -3160 -3500 -3060
rect -3300 -3700 -3200 -3600
rect 4110 -6920 4210 -6820
rect 3680 -10000 3780 -9900
rect 5460 -6320 5560 -6220
rect 20000 -2890 20100 -2790
rect 9150 -8710 9250 -8610
rect 19150 -9100 19250 -9000
rect 19370 -9640 19470 -9540
<< metal3 >>
rect -9600 12399 26800 12400
rect -9600 12340 26805 12399
rect -9600 12300 3780 12340
rect -9600 12100 -9500 12300
rect -9300 12240 3780 12300
rect 3880 12300 26805 12340
rect 3880 12240 26500 12300
rect -9300 12140 26500 12240
rect -9300 12100 3780 12140
rect -9600 12040 3780 12100
rect 3880 12100 26500 12140
rect 26700 12100 26805 12300
rect 3880 12040 26805 12100
rect -9600 12001 26805 12040
rect -9600 12000 26800 12001
rect -8200 10950 25400 11000
rect -8200 10900 14670 10950
rect -8200 10700 -8100 10900
rect -7900 10850 14670 10900
rect 14770 10900 25400 10950
rect 14770 10850 25100 10900
rect -7900 10750 25100 10850
rect -7900 10700 14670 10750
rect -8200 10650 14670 10700
rect 14770 10700 25100 10750
rect 25300 10700 25400 10900
rect 14770 10650 25400 10700
rect -8200 10600 25400 10650
rect -6800 9550 24000 9600
rect -6800 9500 -1330 9550
rect -6800 9300 -6700 9500
rect -6500 9450 -1330 9500
rect -1230 9450 11770 9550
rect 11870 9500 24000 9550
rect 11870 9450 23700 9500
rect -6500 9350 23700 9450
rect -6500 9300 -1330 9350
rect -6800 9250 -1330 9300
rect -1230 9250 11770 9350
rect 11870 9300 23700 9350
rect 23900 9300 24000 9500
rect 11870 9250 24000 9300
rect -6800 9200 24000 9250
rect 11760 8080 11880 8085
rect -1350 8050 -1230 8055
rect -1350 7950 -1340 8050
rect -1240 7950 -1230 8050
rect 11760 7980 11770 8080
rect 11870 7980 11880 8080
rect 11760 7975 11880 7980
rect -1350 7945 -1230 7950
rect -8200 5030 -1180 5080
rect -8200 4930 -8170 5030
rect -8070 4930 -7970 5030
rect -7870 4930 -1330 5030
rect -1230 4930 -1180 5030
rect -8200 4880 -1180 4930
rect 14670 4980 14790 4985
rect 14670 4880 14680 4980
rect 14780 4880 14790 4980
rect 14670 4875 14790 4880
rect 3730 4300 3930 4650
rect 3730 4200 3780 4300
rect 3880 4200 3930 4300
rect 3730 4140 3930 4200
rect 3730 4070 3750 4140
rect 3820 4070 3930 4140
rect 3730 4050 3930 4070
rect 20700 -1350 26800 -1300
rect 20700 -1450 20750 -1350
rect 20850 -1450 26450 -1350
rect 26550 -1450 26650 -1350
rect 26750 -1450 26800 -1350
rect 20700 -1500 26800 -1450
rect 19950 -2790 25400 -2740
rect 19950 -2890 20000 -2790
rect 20100 -2890 25050 -2790
rect 25150 -2890 25250 -2790
rect 25350 -2890 25400 -2790
rect 19950 -2940 25400 -2890
rect -8200 -3060 -3450 -3010
rect -8200 -3160 -8180 -3060
rect -8080 -3160 -7980 -3060
rect -7880 -3160 -3600 -3060
rect -3500 -3160 -3450 -3060
rect -8200 -3210 -3450 -3160
rect -9600 -3600 -3150 -3550
rect -9600 -3610 -3300 -3600
rect -9600 -3710 -9560 -3610
rect -9460 -3710 -9360 -3610
rect -9260 -3700 -3300 -3610
rect -3200 -3700 -3150 -3600
rect -9260 -3710 -3150 -3700
rect -9600 -3750 -3150 -3710
rect 5450 -6220 5570 -6215
rect 5450 -6320 5460 -6220
rect 5560 -6320 5570 -6220
rect 5450 -6325 5570 -6320
rect -9600 -6820 4260 -6770
rect -9600 -6920 -9560 -6820
rect -9460 -6920 -9360 -6820
rect -9260 -6920 4110 -6820
rect 4210 -6920 4260 -6820
rect -9600 -6970 4260 -6920
rect 9140 -8610 9260 -8605
rect 9140 -8710 9150 -8610
rect 9250 -8710 9260 -8610
rect 9140 -8715 9260 -8710
rect 19090 -9000 25400 -8960
rect 19090 -9100 19150 -9000
rect 19250 -9010 25400 -9000
rect 19250 -9100 25050 -9010
rect 19090 -9110 25050 -9100
rect 25150 -9110 25250 -9010
rect 25350 -9110 25400 -9010
rect 19090 -9160 25400 -9110
rect 19320 -9540 26800 -9490
rect 19320 -9640 19370 -9540
rect 19470 -9550 26800 -9540
rect 19470 -9640 26450 -9550
rect 19320 -9650 26450 -9640
rect 26550 -9650 26650 -9550
rect 26750 -9650 26800 -9550
rect 19320 -9690 26800 -9650
rect -8200 -9900 3820 -9850
rect -8200 -10000 -8150 -9900
rect -8050 -10000 -7960 -9900
rect -7860 -10000 3680 -9900
rect 3780 -10000 3820 -9900
rect -8200 -10050 3820 -10000
rect -6800 -14440 24000 -14400
rect -6800 -14500 5460 -14440
rect -6800 -14700 -6700 -14500
rect -6500 -14540 5460 -14500
rect 5560 -14500 24000 -14440
rect 5560 -14540 23700 -14500
rect -6500 -14640 23700 -14540
rect -6500 -14700 5460 -14640
rect -6800 -14740 5460 -14700
rect 5560 -14700 23700 -14640
rect 23900 -14700 24000 -14500
rect 5560 -14740 24000 -14700
rect -6800 -14800 24000 -14740
rect -8200 -15900 25400 -15800
rect -8200 -16100 -8100 -15900
rect -7900 -16100 25100 -15900
rect 25300 -16100 25400 -15900
rect -8200 -16200 25400 -16100
rect -9600 -17230 26800 -17200
rect -9600 -17300 9150 -17230
rect -9600 -17500 -9500 -17300
rect -9300 -17330 9150 -17300
rect 9250 -17300 26800 -17230
rect 9250 -17330 26500 -17300
rect -9300 -17430 26500 -17330
rect -9300 -17500 9150 -17430
rect -9600 -17530 9150 -17500
rect 9250 -17500 26500 -17430
rect 26700 -17500 26800 -17300
rect 9250 -17530 26800 -17500
rect -9600 -17600 26800 -17530
<< via3 >>
rect -9500 12100 -9300 12300
rect 3780 12240 3880 12340
rect 3780 12040 3880 12140
rect 26500 12100 26700 12300
rect -8100 10700 -7900 10900
rect 14670 10850 14770 10950
rect 14670 10650 14770 10750
rect 25100 10700 25300 10900
rect -6700 9300 -6500 9500
rect -1330 9450 -1230 9550
rect 11770 9450 11870 9550
rect -1330 9250 -1230 9350
rect 11770 9250 11870 9350
rect 23700 9300 23900 9500
rect -1340 7950 -1240 8050
rect 11770 7980 11870 8080
rect -8170 4930 -8070 5030
rect -7970 4930 -7870 5030
rect 14680 4880 14780 4980
rect 3780 4200 3880 4300
rect 26450 -1450 26550 -1350
rect 26650 -1450 26750 -1350
rect 25050 -2890 25150 -2790
rect 25250 -2890 25350 -2790
rect -8180 -3160 -8080 -3060
rect -7980 -3160 -7880 -3060
rect -9560 -3710 -9460 -3610
rect -9360 -3710 -9260 -3610
rect 5460 -6320 5560 -6220
rect -9560 -6920 -9460 -6820
rect -9360 -6920 -9260 -6820
rect 9150 -8710 9250 -8610
rect 25050 -9110 25150 -9010
rect 25250 -9110 25350 -9010
rect 26450 -9650 26550 -9550
rect 26650 -9650 26750 -9550
rect -8150 -10000 -8050 -9900
rect -7960 -10000 -7860 -9900
rect -6700 -14700 -6500 -14500
rect 5460 -14540 5560 -14440
rect 5460 -14740 5560 -14640
rect 23700 -14700 23900 -14500
rect -8100 -16100 -7900 -15900
rect 25100 -16100 25300 -15900
rect -9500 -17500 -9300 -17300
rect 9150 -17330 9250 -17230
rect 9150 -17530 9250 -17430
rect 26500 -17500 26700 -17300
<< metal4 >>
rect -9600 12300 -9200 12400
rect -9600 12100 -9500 12300
rect -9300 12100 -9200 12300
rect -9600 -3610 -9200 12100
rect 3730 12340 3930 12400
rect 3730 12240 3780 12340
rect 3880 12240 3930 12340
rect 3730 12140 3930 12240
rect 3730 12040 3780 12140
rect 3880 12040 3930 12140
rect -9600 -3710 -9560 -3610
rect -9460 -3710 -9360 -3610
rect -9260 -3710 -9200 -3610
rect -9600 -6820 -9200 -3710
rect -9600 -6920 -9560 -6820
rect -9460 -6920 -9360 -6820
rect -9260 -6920 -9200 -6820
rect -9600 -17300 -9200 -6920
rect -8200 10900 -7800 11000
rect -8200 10700 -8100 10900
rect -7900 10700 -7800 10900
rect -8200 5030 -7800 10700
rect -8200 4930 -8170 5030
rect -8070 4930 -7970 5030
rect -7870 4930 -7800 5030
rect -8200 -3060 -7800 4930
rect -8200 -3160 -8180 -3060
rect -8080 -3160 -7980 -3060
rect -7880 -3160 -7800 -3060
rect -8200 -9900 -7800 -3160
rect -8200 -10000 -8150 -9900
rect -8050 -10000 -7960 -9900
rect -7860 -10000 -7800 -9900
rect -8200 -15900 -7800 -10000
rect -6800 9500 -6400 9600
rect -6800 9300 -6700 9500
rect -6500 9300 -6400 9500
rect -6800 -14500 -6400 9300
rect -1380 9550 -1180 9600
rect -1380 9450 -1330 9550
rect -1230 9450 -1180 9550
rect -1380 9350 -1180 9450
rect -1380 9250 -1330 9350
rect -1230 9250 -1180 9350
rect -1380 8050 -1180 9250
rect -1380 7950 -1340 8050
rect -1240 7950 -1180 8050
rect -1380 7910 -1180 7950
rect 3730 4300 3930 12040
rect 26400 12300 26800 12400
rect 26400 12100 26500 12300
rect 26700 12100 26800 12300
rect 14620 10950 14820 11000
rect 14620 10850 14670 10950
rect 14770 10850 14820 10950
rect 14620 10750 14820 10850
rect 14620 10650 14670 10750
rect 14770 10650 14820 10750
rect 11720 9550 11920 9600
rect 11720 9450 11770 9550
rect 11870 9450 11920 9550
rect 11720 9350 11920 9450
rect 11720 9250 11770 9350
rect 11870 9250 11920 9350
rect 11720 8080 11920 9250
rect 11720 7980 11770 8080
rect 11870 7980 11920 8080
rect 11720 7910 11920 7980
rect 14620 4980 14820 10650
rect 25000 10900 25400 11000
rect 25000 10700 25100 10900
rect 25300 10700 25400 10900
rect 14620 4880 14680 4980
rect 14780 4880 14820 4980
rect 14620 4830 14820 4880
rect 23600 9500 24000 9600
rect 23600 9300 23700 9500
rect 23900 9300 24000 9500
rect 3730 4200 3780 4300
rect 3880 4200 3930 4300
rect 3730 4050 3930 4200
rect -6800 -14700 -6700 -14500
rect -6500 -14700 -6400 -14500
rect -6800 -14800 -6400 -14700
rect 5410 -6220 5610 -6170
rect 5410 -6320 5460 -6220
rect 5560 -6320 5610 -6220
rect 5410 -14440 5610 -6320
rect 5410 -14540 5460 -14440
rect 5560 -14540 5610 -14440
rect 5410 -14640 5610 -14540
rect 5410 -14740 5460 -14640
rect 5560 -14740 5610 -14640
rect 5410 -14800 5610 -14740
rect 9100 -8610 9300 -8570
rect 9100 -8710 9150 -8610
rect 9250 -8710 9300 -8610
rect -8200 -16100 -8100 -15900
rect -7900 -16100 -7800 -15900
rect -8200 -16200 -7800 -16100
rect -9600 -17500 -9500 -17300
rect -9300 -17500 -9200 -17300
rect -9600 -17600 -9200 -17500
rect 9100 -17230 9300 -8710
rect 23600 -14500 24000 9300
rect 23600 -14700 23700 -14500
rect 23900 -14700 24000 -14500
rect 23600 -14800 24000 -14700
rect 25000 -2790 25400 10700
rect 25000 -2890 25050 -2790
rect 25150 -2890 25250 -2790
rect 25350 -2890 25400 -2790
rect 25000 -9010 25400 -2890
rect 25000 -9110 25050 -9010
rect 25150 -9110 25250 -9010
rect 25350 -9110 25400 -9010
rect 25000 -15900 25400 -9110
rect 25000 -16100 25100 -15900
rect 25300 -16100 25400 -15900
rect 25000 -16200 25400 -16100
rect 26400 -1350 26800 12100
rect 26400 -1450 26450 -1350
rect 26550 -1450 26650 -1350
rect 26750 -1450 26800 -1350
rect 26400 -9550 26800 -1450
rect 26400 -9650 26450 -9550
rect 26550 -9650 26650 -9550
rect 26750 -9650 26800 -9550
rect 9100 -17330 9150 -17230
rect 9250 -17330 9300 -17230
rect 9100 -17430 9300 -17330
rect 9100 -17530 9150 -17430
rect 9250 -17530 9300 -17430
rect 9100 -17600 9300 -17530
rect 26400 -17300 26800 -9650
rect 26400 -17500 26500 -17300
rect 26700 -17500 26800 -17300
rect 26400 -17600 26800 -17500
use count  count_0 ./../count
timestamp 1727161985
transform 1 0 -2340 0 1 -2076
box -880 -3154 3140 -440
use count  count_1
timestamp 1727161985
transform 1 0 16330 0 1 -6486
box -880 -3154 3140 -440
use dco  dco_0 ./../dco
timestamp 1729672293
transform 1 0 2620 0 1 -6850
box 1000 -4280 11940 6160
use qz  qz_0 ./../quantizer
timestamp 1727164310
transform 1 0 15260 0 1 -2230
box 190 -710 5890 730
use vco  vco_0 ./../vco
timestamp 1729655433
transform 1 0 -2020 0 1 680
box 0 0 20640 7330
<< labels >>
rlabel metal2 3480 -7670 3480 -7670 1 D1
rlabel metal2 14720 -9240 14720 -9240 1 p_dco
flabel metal2 20838 7498 21206 8326 1 FreeSans 368 0 0 0 CLK
port 2 nsew signal input
flabel metal2 -3450 7222 -3082 8326 1 FreeSans 368 0 0 0 Anlg_in
port 3 nsew signal input
flabel metal2 -4738 7222 -4370 8326 1 FreeSans 368 0 0 0 ENB
port 5 nsew signal input
flabel metal2 4554 -13570 4830 -13110 1 FreeSans 368 0 0 0 Vbs_12
port 7 nsew signal input
flabel metal2 6486 -13570 6762 -13110 1 FreeSans 368 0 0 0 Vbs_34
port 9 nsew signal input
flabel metal3 -9300 12000 3780 12400 1 FreeSans 736 0 0 0 VCCD
port 4 nsew power input
flabel metal3 -7900 10600 14670 11000 1 FreeSans 736 0 0 0 GND
port 6 nsew ground input
flabel metal3 11870 9200 23700 9600 1 FreeSans 736 0 0 0 VCCA
port 8 nsew power input
flabel metal2 22402 7498 22770 8326 1 FreeSans 368 0 0 0 Dout
port 1 nsew signal output
<< end >>
