* SPICE3 file created from vco.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_po_C4R5Y4 a_n33_165# VSUBS
R0 a_n33_165# a_n33_n595# sky130_fd_pr__res_generic_po w=0.33 l=1.65
.ends

.subckt inv a_0_n1090# a_730_0# a_n80_n1010# w_n120_n40# a_730_n1010# a_n80_0# VSUBS
X0 a_730_n1010# a_0_n1090# a_n80_n1010# VSUBS sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
X1 a_730_0# a_0_n1090# a_n80_0# w_n120_n40# sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
C0 w_n120_n40# VSUBS 3.3756f
.ends

.subckt cc_inv inp inn outp a_2800_1950# a_1840_100# a_n60_1950# a_2800_100# a_n60_100#
+ a_3890_1950# inv_5/VSUBS a_3730_70# a_1840_1950# a_3890_100# w_n60_2030#
Xinv_0 inp inv_1/a_n80_0# a_n60_100# w_n60_2030# inv_1/a_n80_n1010# a_n60_1950# inv_5/VSUBS
+ inv
Xinv_1 inp outp inv_1/a_n80_n1010# w_n60_2030# outp inv_1/a_n80_0# inv_5/VSUBS inv
Xinv_2 outp outp a_1840_100# w_n60_2030# outp a_1840_1950# inv_5/VSUBS inv
Xinv_3 outp outp a_2800_100# w_n60_2030# outp a_2800_1950# inv_5/VSUBS inv
Xinv_4 inn li_4680_1990# a_3890_100# w_n60_2030# inv_5/a_n80_n1010# a_3890_1950# inv_5/VSUBS
+ inv
Xinv_5 inn outp inv_5/a_n80_n1010# w_n60_2030# outp li_4680_1990# inv_5/VSUBS inv
C0 inn outp 2.624074f
C1 inp inv_5/VSUBS 3.826026f
C2 inn inv_5/VSUBS 4.945909f
C3 w_n60_2030# inv_5/VSUBS 19.929615f
C4 outp inv_5/VSUBS 5.266077f
.ends

.subckt ring_osc cc_inv_0/inp cc_inv_4/w_n60_2030# VSUBS
Xcc_inv_0 cc_inv_0/inp cc_inv_0/inp cc_inv_1/inp a_2920_2070# m1_40_n140# a_60_2070#
+ m1_40_n140# m1_40_n140# a_4010_1990# VSUBS cc_inv_0/a_3730_70# a_1960_2070# m1_40_n140#
+ w_60_2070# cc_inv
Xcc_inv_1 cc_inv_1/inp cc_inv_1/inp cc_inv_2/inp cc_inv_1/a_2800_1950# m1_40_n140#
+ cc_inv_1/a_n60_1950# m1_40_n140# m1_40_n140# cc_inv_1/a_3890_1950# VSUBS VSUBS cc_inv_1/a_1840_1950#
+ m1_40_n140# w_60_2070# cc_inv
Xcc_inv_2 cc_inv_2/inp cc_inv_2/inp cc_inv_4/inp cc_inv_2/a_2800_1950# m1_40_n140#
+ cc_inv_2/a_n60_1950# m1_40_n140# m1_40_n140# cc_inv_2/a_3890_1950# VSUBS VSUBS cc_inv_2/a_1840_1950#
+ m1_40_n140# w_60_2070# cc_inv
Xcc_inv_3 cc_inv_3/inp cc_inv_3/inp cc_inv_0/inp cc_inv_3/a_2800_1950# m1_40_n140#
+ cc_inv_3/a_n60_1950# m1_40_n140# m1_40_n140# cc_inv_3/a_3890_1950# VSUBS VSUBS cc_inv_3/a_1840_1950#
+ m1_40_n140# cc_inv_4/w_n60_2030# cc_inv
Xcc_inv_4 cc_inv_4/inp cc_inv_4/inp cc_inv_3/inp cc_inv_4/a_2800_1950# m1_40_n140#
+ cc_inv_4/a_n60_1950# m1_40_n140# m1_40_n140# cc_inv_4/a_3890_1950# VSUBS VSUBS cc_inv_4/a_1840_1950#
+ m1_40_n140# cc_inv_4/w_n60_2030# cc_inv
C0 cc_inv_3/inp VSUBS 13.222344f
C1 cc_inv_4/w_n60_2030# VSUBS 39.86186f
C2 cc_inv_0/inp VSUBS 18.187017f
C3 cc_inv_4/inp VSUBS 17.983839f
C4 cc_inv_2/inp VSUBS 13.158192f
C5 w_60_2070# VSUBS 59.792423f
C6 cc_inv_1/inp VSUBS 13.226386f
C7 m1_40_n140# VSUBS 11.959424f
.ends

.subckt sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
X0 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_204_297# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.149 ps=1.325 w=1 l=0.15
X2 Z A a_204_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3675 ps=1.735 w=1 l=0.15
X3 Z A a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_286_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.23025 ps=1.385 w=0.65 l=0.15
X5 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.23025 pd=1.385 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt vco
Xsky130_fd_pr__res_generic_po_C4R5Y4_0 VSUBS VSUBS sky130_fd_pr__res_generic_po_C4R5Y4
Xsky130_fd_pr__res_generic_po_C4R5Y4_1 VSUBS VSUBS sky130_fd_pr__res_generic_po_C4R5Y4
Xring_osc_0 sky130_fd_sc_hd__einvn_1_0/Z sky130_fd_sc_hd__einvn_1_0/VPB VSUBS ring_osc
Xsky130_fd_sc_hd__einvn_1_0 sky130_fd_sc_hd__einvn_1_0/A sky130_fd_sc_hd__einvn_1_0/TE_B
+ sky130_fd_sc_hd__einvn_1_0/VGND VSUBS sky130_fd_sc_hd__einvn_1_0/VPB sky130_fd_sc_hd__einvn_1_0/VPWR
+ sky130_fd_sc_hd__einvn_1_0/Z sky130_fd_sc_hd__einvn_1
C0 ring_osc_0/cc_inv_3/inp VSUBS 12.886342f
C1 sky130_fd_sc_hd__einvn_1_0/VPB VSUBS 40.348595f
C2 sky130_fd_sc_hd__einvn_1_0/Z VSUBS 17.92247f
C3 ring_osc_0/cc_inv_4/inp VSUBS 17.635897f
C4 ring_osc_0/cc_inv_2/inp VSUBS 12.882699f
C5 ring_osc_0/w_60_2070# VSUBS 59.78896f
C6 ring_osc_0/cc_inv_1/inp VSUBS 12.878458f
C7 ring_osc_0/m1_40_n140# VSUBS 8.633345f
.ends

