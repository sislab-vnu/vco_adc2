magic
tech sky130A
timestamp 1726743291
<< nwell >>
rect 60 1135 125 1295
rect -205 -565 -117 -405
<< pwell >>
rect 40 1015 125 1105
rect -167 -686 -100 -618
<< psubdiff >>
rect 70 1070 100 1085
rect 70 1050 75 1070
rect 95 1050 100 1070
rect 70 1035 100 1050
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
<< nsubdiff >>
rect 70 1195 100 1210
rect 70 1175 75 1195
rect 95 1175 100 1195
rect 70 1160 100 1175
rect -165 -484 -135 -467
rect -165 -501 -158 -484
rect -141 -501 -135 -484
rect -165 -517 -135 -501
<< psubdiffcont >>
rect 75 1050 95 1070
rect -148 -661 -130 -644
<< nsubdiffcont >>
rect 75 1175 95 1195
rect -158 -501 -141 -484
<< locali >>
rect 70 1195 100 1210
rect 70 1175 75 1195
rect 95 1175 100 1195
rect 70 1160 100 1175
rect -10 1114 135 1135
rect 70 1070 100 1085
rect 70 1050 75 1070
rect 95 1050 100 1070
rect 70 1035 100 1050
rect -165 -484 -135 -467
rect 120 -480 175 -450
rect -165 -501 -158 -484
rect -141 -501 -135 -484
rect -165 -517 -135 -501
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
<< viali >>
rect 75 1175 95 1195
rect -122 1112 -105 1129
rect 75 1050 95 1070
rect -70 -590 -50 -570
rect 99 -589 116 -572
rect -148 -661 -130 -644
<< metal1 >>
rect 70 1195 100 1210
rect 70 1175 75 1195
rect 95 1175 100 1195
rect 70 1160 100 1175
rect -165 1129 -97 1139
rect -165 1112 -122 1129
rect -105 1112 -97 1129
rect -165 1103 -97 1112
rect 70 1070 100 1085
rect 70 1050 75 1070
rect 95 1050 100 1070
rect 70 1035 100 1050
rect -165 -517 -135 -467
rect -90 -570 -47 -555
rect -140 -590 -70 -570
rect -50 -590 -47 -570
rect -140 -600 -47 -590
rect 96 -571 121 -558
rect 96 -572 165 -571
rect 96 -589 99 -572
rect 116 -589 165 -572
rect 96 -605 121 -589
rect -156 -644 -125 -627
rect -156 -661 -148 -644
rect -130 -661 -125 -644
rect -156 -677 -125 -661
use dco_freq  dco_freq_0
timestamp 1726743291
transform 1 0 4160 0 1 25
box -440 -625 1665 320
use dco_freq  dco_freq_1
timestamp 1726743291
transform 1 0 4160 0 1 -1145
box -440 -625 1665 320
use dco_idac  dco_idac_0
timestamp 1726728476
transform 1 0 1430 0 1 -30
box -930 -1580 1610 370
use dco_ring_osc  dco_ring_osc_0
timestamp 1726107115
transform 1 0 840 0 1 2003
box -250 -1260 4720 1080
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -141 0 1 1004
box -19 -24 203 296
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -101 0 1 -696
box -19 -24 249 296
<< end >>
