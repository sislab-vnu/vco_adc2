** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/DLib_UpDownCounter.sch
.subckt DLib_UpDownCounter UP DOWN setB Dout_buf VDDA GND
*.PININFO DOWN:I Dout_buf:O GND:I setB:I UP:I VDDA:I
X_inv_0 setB GND GND VDDA VDDA setBi sky130_fd_sc_hd__inv_2
X_upFF UP_buf Q2N setBi GND GND VDDA VDDA Q1 sky130_fd_sc_hd__dfstp_1
X_dwFF DWN_buf Q1_buf setBi GND GND VDDA VDDA Q2 sky130_fd_sc_hd__dfstp_1
x5 Q1 Q2 GND GND VDDA VDDA Dout sky130_fd_sc_hd__xor2_1
X_buf_3 UP GND GND VDDA VDDA UP_buf sky130_fd_sc_hd__buf_2
X_buf_4 Q1 GND GND VDDA VDDA Q1_buf sky130_fd_sc_hd__buf_2
X_buf_5 Dout GND GND VDDA VDDA Dout_buf sky130_fd_sc_hd__buf_2
X_buf_6 DOWN GND GND VDDA VDDA DWN_buf sky130_fd_sc_hd__buf_2
X_inv_1 Q2 GND GND VDDA VDDA Q2N sky130_fd_sc_hd__inv_2
.ends
.end
