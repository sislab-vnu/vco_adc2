** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/DLib_UpDownCounter_tb.sch
**.subckt DLib_UpDownCounter_tb
x2 UP Anlg_in ENB VDDA GND ALib_VCO
x1 VDDA GND UP ENB DOWN Dout DLib_UpDownCounter
V1 Anlg_in GND DC=0 sin(0.8 0.4 0.5Meg 0 0 0)
V2 VDDA GND DC=1.8
V3 ENB GND DC=0 PULSE(0 1.8 0 0.1n 0.1n 20n 1)
V4 DOWN GND DC=0 PULSE(0 1.8 0 0.1n 0.1n 17n 41.67n)
**** begin user architecture code


.lib /home/dkits/openpdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /home/dkits/openpdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice




.control
set num_threads=10
save all
TRAN 1n 10u
.endc


**** end user architecture code
**.ends

* expanding   symbol:  ALib_VCO.sym # of pins=5
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/ALib_VCO.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/ALib_VCO.sch
.subckt ALib_VCO p[4] Anlg_in ENB VDDA GND
*.ipin Anlg_in
*.ipin VDDA
*.ipin ENB
*.opin p[4]
*.ipin GND
Xro_1 net1 VDDA p[0] p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4] GND 5s_cc_osc
x1 VDDA ENB VGND VNB VPB VPWR pn[4] sky130_fd_sc_hd__einvp_1
R1 net1 Anlg_in sky130_fd_pr__res_generic_po W=1 L=1 m=1
R2 net2 net1 sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends


* expanding   symbol:  DLib_UpDownCounter.sym # of pins=6
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/DLib_UpDownCounter.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/DLib_UpDownCounter.sch
.subckt DLib_UpDownCounter VDDA GND UP setB DOWN Dout_buf
*.ipin DOWN
*.opin Dout_buf
*.ipin GND
*.ipin setB
*.ipin UP
*.ipin VDDA
X_inv_0 setB GND GND VDDA VDDA setBi sky130_fd_sc_hd__inv_2
X_upFF UP_buf Q2N setBi GND GND VDDA VDDA Q1 sky130_fd_sc_hd__dfstp_1
X_dwFF DWN_buf Q1_buf setBi GND GND VDDA VDDA Q2 sky130_fd_sc_hd__dfstp_1
x5 Q1 Q2 GND GND VDDA VDDA Dout sky130_fd_sc_hd__xor2_1
X_buf_3 UP GND GND VDDA VDDA UP_buf sky130_fd_sc_hd__buf_2
X_buf_4 Q1 GND GND VDDA VDDA Q1_buf sky130_fd_sc_hd__buf_2
X_buf_5 Dout GND GND VDDA VDDA Dout_buf sky130_fd_sc_hd__buf_2
X_buf_6 DOWN GND GND VDDA VDDA DWN_buf sky130_fd_sc_hd__buf_2
X_inv_1 Q2 GND GND VDDA VDDA Q2N sky130_fd_sc_hd__inv_2
.ends


* expanding   symbol:  5s_cc_osc.sym # of pins=13
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/5s_cc_osc.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/5s_cc_osc.sch
.subckt 5s_cc_osc VGND VDDA p[0] p[1] p[2] p[3] p[4] pn[0] pn[1] pn[2] pn[3] pn[4] GND
*.iopin VDDA
*.iopin VGND
*.opin pn[0]
*.iopin p[0]
*.opin pn[1]
*.opin p[1]
*.opin p[2]
*.opin p[3]
*.opin p[4]
*.opin pn[2]
*.opin pn[3]
*.opin pn[4]
*.iopin GND
Xi_1 p[4] pn[4] VDDA VGND p[0] pn[0] GND cc_inv
Xi_2 p[0] pn[0] VDDA VGND p[1] pn[1] GND cc_inv
Xi_3 p[1] pn[1] VDDA VGND p[2] pn[2] GND cc_inv
Xi_4 p[2] pn[2] VDDA VGND p[3] pn[3] GND cc_inv
Xi_6 p[3] pn[3] VDDA VGND p[4] pn[4] GND cc_inv
.ends


* expanding   symbol:  cc_inv.sym # of pins=7
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/cc_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/cc_inv.sch
.subckt cc_inv inp inn VDDA VGND outp outn GND
*.opin outp
*.ipin inn
*.iopin VGND
*.opin outn
*.ipin inp
*.iopin VDDA
*.iopin GND
Xi_1 VDDA VGND outp GND inp main_inv
Xi_2 VDDA VGND outn GND inn main_inv
Xi_3 VDDA VGND outn GND outp aux_inv
Xi_4 VDDA VGND outp GND outn aux_inv
.ends


* expanding   symbol:  main_inv.sym # of pins=5
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/main_inv.sch
.subckt main_inv VDDA VGND Y GND A
*.iopin VDDA
*.iopin VGND
*.ipin A
*.opin Y
*.iopin GND
XM1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  aux_inv.sym # of pins=5
** sym_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sym
** sch_path: /home/userdata/k63D/toind_63d/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sch
.subckt aux_inv VDDA VGND Y GND A
*.iopin VDDA
*.iopin VGND
*.ipin A
*.opin Y
*.iopin GND
XM1 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
