** sch_path: /home/toind/work/sislab_vnu/vco_adc2/xschem/lib/aux_inv.sch
.subckt aux_inv A Y VGND VDDA GND
*.PININFO VDDA:B VGND:B A:I Y:O GND:B
XM3 Y A VGND GND sky130_fd_pr__nfet_01v8 L=3.65 W=4 nf=1 m=1
XM2 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=3.65 W=5 nf=1 m=1
.ends
.end
