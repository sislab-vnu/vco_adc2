* this file contains all analog circuits written by SPICE
* lib 	: analog_library
* tech	: 130nm Skywater
* author: Duc-Manh Tran

* Subcircuit    : inv_12
*****************************************************************************
.subckt inv_12 y a VDDPIN  VSSPIN VNBPIN
XM1 a y VSSPIN VNBPIN sky130_fd_pr__nfet_01v8 w=4.5 l=1.8 nf=4
XM2 a y VDDPIN VDDPIN sky130_fd_pr__pfet_01v8 w=4.5 l=1.8 nf=2
.ends

* Subcircuit    : inv_34
*****************************************************************************
.subckt inv_34 y a VDDPIN  VSSPIN VNBPIN
XM1 a y VSSPIN VNBPIN sky130_fd_pr__nfet_01v8 w=4 l=1.8 nf=2
XM2 a y VDDPIN VDDPIN sky130_fd_pr__pfet_01v8 w=4 l=1.8 nf=1
.ends

* Subcircuit    : cc_inv
*******************************************************************************
.subckt cc_inv inp inn outp outn vdd vss VSUBS
xi1 inp outp vdd vss VSUBS inv_12
xi2 inn outn vdd vss VSUBS inv_12
xi3 outp outn vdd vss VSUBS inv_34
xi4 outn outp vdd vss VSUBS inv_34
.ends

* Subcircuit    : ring_osc
********************************************************************************
.subckt ring_osc p[0] p[1] p[2] p[3] p[4] input enb vdd VSUBS
Xc2 p[0] p_n[0] p[1] p_n[1] vdd input VSUBS cc_inv
Xc3 p[1] p_n[1] p[2] p_n[2] vdd input VSUBS cc_inv
Xc4 p[2] p_n[2] p[3] p_n[3] vdd input VSUBS cc_inv
Xc5 p[3] p_n[3] p[4] p_n[4] vdd input VSUBS cc_inv
Xc6 p[4] p_n[4] p[0] p_n[0] vdd input VSUBS cc_inv
.ends

.subckt vco p[0] p[1] p[2] p[3] p[4] input enb vdd vss v_ctr
Xro_1 p[0] p[1] p[2] p[3] p[4] vdd vss v_ctr ring_osc
Xconb_1 vss VSUBS vdd vdd hi_logic lo_logic sky130_fd_sc_hd__conb_1
Xeinvp_1 hi_logic enb vss VSUBS vdd vdd p[0] sky130_fd_sc_hd__einvp_1
R0 v_ctr input sky130_fd_pr__res_generic_po w=2e+06u l=4.15e+06u
R1 v_ctr vss sky130_fd_pr__res_generic_po w=2e+06u l=4.15e+06u
.ends

