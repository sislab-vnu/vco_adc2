VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO count
  CLASS BLOCK ;
  FOREIGN count ;
  ORIGIN 4.400 15.770 ;
  SIZE 20.100 BY 13.570 ;
  PIN UP
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT -4.400 -4.150 -3.050 -3.800 ;
        RECT -3.425 -4.175 -3.070 -4.150 ;
    END
  END UP
  PIN SetB
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT -3.255 -9.295 -2.925 -9.045 ;
      LAYER met1 ;
        RECT -4.150 -9.350 -2.900 -9.000 ;
    END
  END SetB
  PIN DOWN
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 13.600 -13.790 14.150 -13.750 ;
        RECT 12.960 -14.170 14.150 -13.790 ;
        RECT 13.600 -14.200 14.150 -14.170 ;
    END
  END DOWN
  PIN Dout_buf
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 10.290 -9.280 10.545 -8.375 ;
        RECT 10.375 -10.010 10.545 -9.280 ;
        RECT 10.290 -10.585 10.545 -10.010 ;
      LAYER met1 ;
        RECT 10.250 -9.450 10.550 -8.750 ;
        RECT 10.250 -9.800 11.400 -9.450 ;
        RECT 10.250 -9.810 10.550 -9.800 ;
    END
  END Dout_buf
  PIN GND
    ANTENNADIFFAREA 5.467100 ;
    PORT
      LAYER pwell ;
        RECT -3.020 -4.350 -1.675 -4.145 ;
        RECT -4.300 -4.375 -3.450 -4.350 ;
        RECT -3.020 -4.375 -0.050 -4.350 ;
        RECT 1.295 -4.375 2.215 -4.155 ;
        RECT 8.295 -4.255 9.215 -4.145 ;
        RECT 6.880 -4.350 9.215 -4.255 ;
        RECT 6.880 -4.375 11.450 -4.350 ;
        RECT 11.890 -4.375 13.235 -4.145 ;
        RECT -4.300 -5.050 13.235 -4.375 ;
        RECT -3.505 -5.055 -1.675 -5.050 ;
        RECT -0.065 -5.055 9.215 -5.050 ;
        RECT 11.405 -5.055 13.235 -5.050 ;
        RECT -3.365 -5.245 -3.195 -5.055 ;
        RECT 0.075 -5.245 0.245 -5.055 ;
        RECT 11.545 -5.245 11.715 -5.055 ;
        RECT -4.250 -9.355 -3.300 -9.350 ;
        RECT -4.250 -10.250 -1.995 -9.355 ;
        RECT -3.345 -10.265 -1.995 -10.250 ;
        RECT 4.695 -10.050 7.865 -9.825 ;
        RECT 4.695 -10.055 9.250 -10.050 ;
        RECT 9.720 -10.055 11.065 -9.825 ;
        RECT -3.215 -10.455 -3.045 -10.265 ;
        RECT 4.695 -10.735 11.065 -10.055 ;
        RECT 4.795 -10.925 4.965 -10.735 ;
        RECT 7.850 -10.750 9.250 -10.735 ;
        RECT 9.375 -10.925 9.545 -10.735 ;
        RECT -1.435 -12.915 -1.265 -12.725 ;
        RECT -1.150 -12.915 0.350 -12.900 ;
        RECT 9.315 -12.915 9.485 -12.725 ;
        RECT 9.600 -12.915 11.600 -12.900 ;
        RECT 13.085 -12.915 13.255 -12.725 ;
        RECT -2.485 -13.595 13.395 -12.915 ;
        RECT -2.485 -13.715 2.680 -13.595 ;
        RECT -2.485 -13.825 1.265 -13.715 ;
        RECT 7.345 -13.815 8.265 -13.595 ;
        RECT 9.600 -13.600 12.910 -13.595 ;
        RECT 11.565 -13.825 12.910 -13.600 ;
        RECT -1.150 -13.850 0.350 -13.825 ;
      LAYER li1 ;
        RECT -4.100 -4.900 -3.700 -4.400 ;
        RECT -2.950 -5.075 -2.620 -4.695 ;
        RECT -2.020 -4.900 -1.760 -4.235 ;
        RECT -2.020 -5.075 -0.050 -4.900 ;
        RECT 0.445 -5.075 0.775 -4.695 ;
        RECT 1.385 -5.075 1.715 -4.695 ;
        RECT 3.540 -5.075 3.950 -4.635 ;
        RECT 4.690 -5.075 5.010 -4.615 ;
        RECT 6.620 -5.075 7.280 -4.595 ;
        RECT 8.410 -5.075 8.695 -4.615 ;
        RECT 9.550 -5.075 11.400 -4.950 ;
        RECT 11.960 -5.075 12.290 -4.695 ;
        RECT 12.890 -5.075 13.150 -4.235 ;
        RECT -3.510 -5.245 13.240 -5.075 ;
        RECT -1.800 -5.400 -0.050 -5.245 ;
        RECT 9.550 -5.400 11.400 -5.245 ;
        RECT -4.050 -10.100 -3.650 -9.600 ;
        RECT -3.235 -10.285 -3.005 -9.465 ;
        RECT -2.335 -10.100 -2.125 -9.465 ;
        RECT -2.335 -10.285 2.550 -10.100 ;
        RECT -3.360 -10.450 2.550 -10.285 ;
        RECT -3.360 -10.455 -1.980 -10.450 ;
        RECT 2.200 -10.650 2.550 -10.450 ;
        RECT 4.785 -10.650 5.115 -10.365 ;
        RECT 2.200 -10.755 5.115 -10.650 ;
        RECT 5.625 -10.755 5.955 -10.365 ;
        RECT 7.495 -10.755 7.785 -9.920 ;
        RECT 8.300 -10.600 8.800 -10.200 ;
        RECT 9.790 -10.755 10.120 -10.375 ;
        RECT 10.720 -10.755 10.980 -9.915 ;
        RECT 2.200 -10.925 7.870 -10.755 ;
        RECT 9.230 -10.925 11.070 -10.755 ;
        RECT 2.200 -11.000 4.850 -10.925 ;
        RECT -1.250 -12.725 0.050 -12.600 ;
        RECT 2.200 -12.725 2.550 -11.000 ;
        RECT 9.600 -12.725 11.750 -12.700 ;
        RECT -2.500 -12.895 13.400 -12.725 ;
        RECT -2.355 -13.715 -2.145 -12.895 ;
        RECT -1.475 -13.050 0.050 -12.895 ;
        RECT -1.475 -13.715 -1.245 -13.050 ;
        RECT 0.865 -13.355 1.150 -12.895 ;
        RECT 2.280 -13.375 2.940 -12.895 ;
        RECT 4.550 -13.355 4.870 -12.895 ;
        RECT 5.610 -13.335 6.020 -12.895 ;
        RECT 7.845 -13.275 8.175 -12.895 ;
        RECT 8.785 -13.275 9.115 -12.895 ;
        RECT 9.600 -13.050 11.910 -12.895 ;
        RECT 10.700 -13.450 11.200 -13.050 ;
        RECT 11.650 -13.735 11.910 -13.050 ;
        RECT 12.510 -13.275 12.840 -12.895 ;
      LAYER met1 ;
        RECT -4.100 -4.900 -3.700 -4.400 ;
        RECT -4.100 -4.920 -3.400 -4.900 ;
        RECT -4.100 -5.400 -1.670 -4.920 ;
        RECT -0.070 -5.400 9.590 -4.920 ;
        RECT 11.400 -5.400 13.240 -4.920 ;
        RECT -4.050 -10.100 -3.650 -9.600 ;
        RECT -4.050 -10.130 -3.350 -10.100 ;
        RECT -4.050 -10.610 -1.980 -10.130 ;
        RECT 2.200 -10.450 2.550 -5.400 ;
        RECT 8.300 -10.600 8.800 -10.200 ;
        RECT -4.050 -10.650 -3.350 -10.610 ;
        RECT 4.650 -11.080 11.070 -10.600 ;
        RECT 7.850 -11.100 9.250 -11.080 ;
        RECT -2.500 -13.050 -1.120 -12.570 ;
        RECT -0.030 -13.050 9.630 -12.570 ;
        RECT 11.560 -13.050 13.400 -12.570 ;
        RECT 10.700 -13.450 11.200 -13.050 ;
    END
  END GND
  PIN VCCD
    ANTENNADIFFAREA 7.256200 ;
    PORT
      LAYER nwell ;
        RECT -4.300 -3.900 13.450 -2.200 ;
        RECT -4.250 -7.460 -3.350 -7.400 ;
        RECT -4.250 -9.065 -1.790 -7.460 ;
        RECT 8.050 -7.930 9.050 -7.900 ;
        RECT -4.250 -9.100 -3.400 -9.065 ;
        RECT 4.460 -9.535 11.260 -7.930 ;
        RECT 8.050 -9.550 9.050 -9.535 ;
        RECT -0.950 -14.115 -0.100 -14.100 ;
        RECT 9.800 -14.115 11.600 -14.100 ;
        RECT -2.690 -15.720 13.590 -14.115 ;
        RECT -0.950 -15.750 -0.100 -15.720 ;
        RECT 9.800 -15.750 11.750 -15.720 ;
      LAYER li1 ;
        RECT 13.150 -2.355 15.700 -2.350 ;
        RECT -3.510 -2.525 -1.670 -2.355 ;
        RECT -0.070 -2.525 9.590 -2.355 ;
        RECT 11.400 -2.525 15.700 -2.355 ;
        RECT -2.950 -3.285 -2.620 -2.525 ;
        RECT -2.020 -3.675 -1.760 -2.525 ;
        RECT -1.050 -3.300 -0.650 -2.800 ;
        RECT 0.445 -3.025 0.775 -2.525 ;
        RECT 1.385 -3.025 1.715 -2.525 ;
        RECT 3.360 -2.905 3.740 -2.525 ;
        RECT 4.260 -2.905 4.590 -2.525 ;
        RECT 5.870 -2.905 6.290 -2.525 ;
        RECT 6.960 -3.215 7.290 -2.525 ;
        RECT 8.410 -3.325 8.695 -2.525 ;
        RECT 11.960 -3.285 12.290 -2.525 ;
        RECT 12.890 -2.700 15.700 -2.525 ;
        RECT 12.890 -3.675 13.150 -2.700 ;
        RECT -2.150 -7.565 5.000 -7.550 ;
        RECT -3.360 -7.735 5.000 -7.565 ;
        RECT -4.050 -8.350 -3.650 -7.850 ;
        RECT -3.235 -8.875 -3.005 -7.735 ;
        RECT -2.335 -7.900 5.000 -7.735 ;
        RECT -2.335 -8.875 -2.125 -7.900 ;
        RECT 4.650 -8.035 5.000 -7.900 ;
        RECT 4.650 -8.205 7.870 -8.035 ;
        RECT 9.230 -8.050 11.070 -8.035 ;
        RECT 15.350 -8.050 15.700 -2.700 ;
        RECT 9.230 -8.205 15.700 -8.050 ;
        RECT 5.705 -9.055 5.875 -8.205 ;
        RECT 6.545 -8.715 6.715 -8.205 ;
        RECT 8.400 -9.100 8.800 -8.600 ;
        RECT 9.790 -8.965 10.120 -8.205 ;
        RECT 10.720 -8.400 15.700 -8.205 ;
        RECT 10.720 -9.355 10.980 -8.400 ;
        RECT -2.355 -15.445 -2.145 -14.305 ;
        RECT -1.475 -15.445 -1.245 -14.305 ;
        RECT -0.650 -15.050 -0.250 -14.550 ;
        RECT 0.865 -15.445 1.150 -14.645 ;
        RECT 2.270 -15.445 2.600 -14.755 ;
        RECT 3.270 -15.445 3.690 -15.065 ;
        RECT 4.970 -15.445 5.300 -15.065 ;
        RECT 5.820 -15.445 6.200 -15.065 ;
        RECT 7.845 -15.445 8.175 -14.945 ;
        RECT 8.785 -15.445 9.115 -14.945 ;
        RECT 11.650 -15.445 11.910 -14.295 ;
        RECT 12.510 -15.445 12.840 -14.685 ;
        RECT 15.350 -15.400 15.700 -8.400 ;
        RECT 13.350 -15.445 15.700 -15.400 ;
        RECT -2.500 -15.615 -1.120 -15.445 ;
        RECT -0.030 -15.615 9.630 -15.445 ;
        RECT 11.560 -15.615 15.700 -15.445 ;
        RECT 13.350 -15.750 15.700 -15.615 ;
      LAYER met1 ;
        RECT -3.510 -2.680 13.240 -2.200 ;
        RECT -1.700 -2.700 0.000 -2.680 ;
        RECT 9.550 -2.700 11.400 -2.680 ;
        RECT -1.050 -3.300 -0.650 -2.700 ;
        RECT -4.050 -7.410 -3.300 -7.400 ;
        RECT -4.050 -7.890 -1.980 -7.410 ;
        RECT 7.850 -7.880 9.250 -7.850 ;
        RECT -4.050 -7.900 -3.300 -7.890 ;
        RECT -4.050 -8.350 -3.650 -7.900 ;
        RECT 4.650 -8.350 11.070 -7.880 ;
        RECT 4.650 -8.360 7.870 -8.350 ;
        RECT 8.400 -9.100 8.800 -8.350 ;
        RECT 9.230 -8.360 11.070 -8.350 ;
        RECT -2.500 -15.300 -1.120 -15.290 ;
        RECT -0.650 -15.300 -0.250 -14.550 ;
        RECT -0.030 -15.300 9.630 -15.290 ;
        RECT 11.560 -15.300 13.400 -15.290 ;
        RECT -2.500 -15.750 13.400 -15.300 ;
        RECT -2.500 -15.770 -1.120 -15.750 ;
        RECT -0.030 -15.770 9.630 -15.750 ;
        RECT 11.560 -15.770 13.400 -15.750 ;
    END
  END VCCD
  OBS
      LAYER li1 ;
        RECT -3.335 -3.455 -3.165 -2.695 ;
        RECT -3.335 -3.625 -2.620 -3.455 ;
        RECT -2.450 -3.600 -2.195 -2.695 ;
        RECT 0.105 -3.195 0.275 -2.695 ;
        RECT 0.105 -3.365 0.770 -3.195 ;
        RECT -2.790 -3.835 -2.620 -3.625 ;
        RECT -2.790 -4.165 -2.535 -3.835 ;
        RECT -2.365 -3.850 -2.195 -3.600 ;
        RECT 0.020 -3.850 0.370 -3.535 ;
        RECT -2.365 -4.050 0.370 -3.850 ;
        RECT -2.790 -4.355 -2.620 -4.165 ;
        RECT -2.365 -4.330 -2.195 -4.050 ;
        RECT 0.020 -4.185 0.370 -4.050 ;
        RECT -3.335 -4.525 -2.620 -4.355 ;
        RECT -3.335 -4.905 -3.165 -4.525 ;
        RECT -2.450 -4.905 -2.195 -4.330 ;
        RECT 0.540 -4.355 0.770 -3.365 ;
        RECT 0.105 -4.525 0.770 -4.355 ;
        RECT 0.105 -4.815 0.275 -4.525 ;
        RECT 0.945 -4.815 1.170 -2.695 ;
        RECT 1.885 -3.195 2.055 -2.695 ;
        RECT 2.290 -2.910 3.120 -2.740 ;
        RECT 1.360 -3.365 2.055 -3.195 ;
        RECT 1.360 -4.335 1.530 -3.365 ;
        RECT 1.700 -4.155 2.110 -3.535 ;
        RECT 2.280 -3.585 2.780 -3.205 ;
        RECT 1.360 -4.525 2.055 -4.335 ;
        RECT 2.280 -4.455 2.500 -3.585 ;
        RECT 2.950 -3.755 3.120 -2.910 ;
        RECT 3.920 -3.075 4.090 -2.785 ;
        RECT 5.060 -2.995 5.690 -2.745 ;
        RECT 5.520 -3.075 5.690 -2.995 ;
        RECT 6.490 -3.075 6.730 -2.785 ;
        RECT 3.290 -3.325 4.660 -3.075 ;
        RECT 3.290 -3.585 3.540 -3.325 ;
        RECT 4.050 -3.755 4.300 -3.595 ;
        RECT 2.950 -3.925 4.300 -3.755 ;
        RECT 2.950 -3.965 3.370 -3.925 ;
        RECT 2.680 -4.515 3.030 -4.145 ;
        RECT 1.885 -4.855 2.055 -4.525 ;
        RECT 3.200 -4.695 3.370 -3.965 ;
        RECT 4.470 -4.095 4.660 -3.325 ;
        RECT 3.540 -4.425 3.950 -4.095 ;
        RECT 2.355 -4.895 3.370 -4.695 ;
        RECT 4.240 -4.435 4.660 -4.095 ;
        RECT 4.830 -3.505 5.350 -3.195 ;
        RECT 5.520 -3.245 6.730 -3.075 ;
        RECT 4.830 -4.265 5.000 -3.505 ;
        RECT 5.170 -4.095 5.350 -3.685 ;
        RECT 5.520 -3.755 5.690 -3.245 ;
        RECT 7.460 -3.395 7.630 -2.785 ;
        RECT 7.900 -3.245 8.230 -2.735 ;
        RECT 7.460 -3.415 7.780 -3.395 ;
        RECT 5.860 -3.585 7.780 -3.415 ;
        RECT 5.520 -3.925 7.420 -3.755 ;
        RECT 5.750 -4.265 6.080 -4.145 ;
        RECT 4.830 -4.435 6.080 -4.265 ;
        RECT 4.240 -4.865 4.490 -4.435 ;
        RECT 6.250 -4.685 6.420 -3.925 ;
        RECT 7.090 -3.985 7.420 -3.925 ;
        RECT 6.610 -4.155 6.940 -4.095 ;
        RECT 6.610 -4.425 7.270 -4.155 ;
        RECT 7.590 -4.480 7.780 -3.585 ;
        RECT 5.570 -4.855 6.420 -4.685 ;
        RECT 7.460 -4.810 7.780 -4.480 ;
        RECT 7.980 -3.835 8.230 -3.245 ;
        RECT 8.875 -3.505 9.130 -2.835 ;
        RECT 8.950 -3.800 9.130 -3.505 ;
        RECT 11.575 -3.455 11.745 -2.695 ;
        RECT 11.575 -3.625 12.290 -3.455 ;
        RECT 12.460 -3.600 12.715 -2.695 ;
        RECT 8.950 -3.805 11.500 -3.800 ;
        RECT 7.980 -4.165 8.780 -3.835 ;
        RECT 7.980 -4.815 8.230 -4.165 ;
        RECT 8.950 -4.175 11.840 -3.805 ;
        RECT 12.120 -3.835 12.290 -3.625 ;
        RECT 12.120 -4.165 12.375 -3.835 ;
        RECT 8.950 -4.200 11.500 -4.175 ;
        RECT 8.950 -4.365 9.130 -4.200 ;
        RECT 12.120 -4.355 12.290 -4.165 ;
        RECT 12.545 -4.330 12.715 -3.600 ;
        RECT 8.875 -4.895 9.130 -4.365 ;
        RECT 11.575 -4.525 12.290 -4.355 ;
        RECT 11.575 -4.905 11.745 -4.525 ;
        RECT 12.460 -4.905 12.715 -4.330 ;
        RECT -2.835 -8.885 -2.505 -7.905 ;
        RECT -2.755 -9.100 -2.505 -8.885 ;
        RECT 4.735 -9.055 5.115 -8.375 ;
        RECT 6.045 -8.885 6.375 -8.375 ;
        RECT 6.885 -8.885 7.285 -8.375 ;
        RECT 6.045 -9.055 7.285 -8.885 ;
        RECT -2.755 -9.270 -2.500 -9.100 ;
        RECT -2.755 -9.485 -2.505 -9.270 ;
        RECT -2.835 -10.115 -2.505 -9.485 ;
        RECT 4.735 -10.015 4.905 -9.055 ;
        RECT 5.075 -9.395 6.380 -9.225 ;
        RECT 7.465 -9.305 7.785 -8.375 ;
        RECT 9.405 -9.135 9.575 -8.375 ;
        RECT 9.405 -9.305 10.120 -9.135 ;
        RECT 5.075 -9.845 5.320 -9.395 ;
        RECT 5.490 -9.765 6.040 -9.565 ;
        RECT 6.210 -9.595 6.380 -9.395 ;
        RECT 7.155 -9.450 7.785 -9.305 ;
        RECT 7.155 -9.500 9.000 -9.450 ;
        RECT 9.315 -9.500 9.670 -9.485 ;
        RECT 6.210 -9.765 6.585 -9.595 ;
        RECT 6.755 -10.015 6.985 -9.515 ;
        RECT 4.735 -10.185 6.985 -10.015 ;
        RECT 7.155 -9.700 9.670 -9.500 ;
        RECT 5.285 -10.505 5.455 -10.185 ;
        RECT 7.155 -10.355 7.325 -9.700 ;
        RECT 9.315 -9.855 9.670 -9.700 ;
        RECT 9.950 -9.515 10.120 -9.305 ;
        RECT 9.950 -9.845 10.205 -9.515 ;
        RECT 9.950 -10.035 10.120 -9.845 ;
        RECT 6.370 -10.525 7.325 -10.355 ;
        RECT 9.405 -10.205 10.120 -10.035 ;
        RECT 9.405 -10.585 9.575 -10.205 ;
        RECT -1.975 -13.695 -1.645 -13.065 ;
        RECT 0.430 -13.605 0.685 -13.075 ;
        RECT -1.975 -14.295 -1.725 -13.695 ;
        RECT -1.555 -13.890 -1.225 -13.885 ;
        RECT 0.430 -13.890 0.610 -13.605 ;
        RECT 1.330 -13.805 1.580 -13.155 ;
        RECT -1.555 -14.130 0.610 -13.890 ;
        RECT -1.555 -14.135 -1.225 -14.130 ;
        RECT -1.975 -15.275 -1.645 -14.295 ;
        RECT 0.430 -14.465 0.610 -14.130 ;
        RECT 0.780 -14.135 1.580 -13.805 ;
        RECT 0.430 -15.135 0.685 -14.465 ;
        RECT 1.330 -14.725 1.580 -14.135 ;
        RECT 1.780 -13.490 2.100 -13.160 ;
        RECT 3.140 -13.285 3.990 -13.115 ;
        RECT 1.780 -14.385 1.970 -13.490 ;
        RECT 2.290 -13.815 2.950 -13.545 ;
        RECT 2.620 -13.875 2.950 -13.815 ;
        RECT 2.140 -14.045 2.470 -13.985 ;
        RECT 3.140 -14.045 3.310 -13.285 ;
        RECT 5.070 -13.535 5.320 -13.105 ;
        RECT 3.480 -13.705 4.730 -13.535 ;
        RECT 3.480 -13.825 3.810 -13.705 ;
        RECT 2.140 -14.215 4.040 -14.045 ;
        RECT 1.780 -14.555 3.700 -14.385 ;
        RECT 1.780 -14.575 2.100 -14.555 ;
        RECT 1.330 -15.235 1.660 -14.725 ;
        RECT 1.930 -15.185 2.100 -14.575 ;
        RECT 3.870 -14.725 4.040 -14.215 ;
        RECT 4.210 -14.285 4.390 -13.875 ;
        RECT 4.560 -14.465 4.730 -13.705 ;
        RECT 2.830 -14.895 4.040 -14.725 ;
        RECT 4.210 -14.775 4.730 -14.465 ;
        RECT 4.900 -13.875 5.320 -13.535 ;
        RECT 6.190 -13.275 7.205 -13.075 ;
        RECT 5.610 -13.875 6.020 -13.545 ;
        RECT 4.900 -14.645 5.090 -13.875 ;
        RECT 6.190 -14.005 6.360 -13.275 ;
        RECT 7.505 -13.445 7.675 -13.115 ;
        RECT 6.530 -13.825 6.880 -13.455 ;
        RECT 6.190 -14.045 6.610 -14.005 ;
        RECT 5.260 -14.215 6.610 -14.045 ;
        RECT 5.260 -14.375 5.510 -14.215 ;
        RECT 6.020 -14.645 6.270 -14.385 ;
        RECT 4.900 -14.895 6.270 -14.645 ;
        RECT 2.830 -15.185 3.070 -14.895 ;
        RECT 3.870 -14.975 4.040 -14.895 ;
        RECT 3.870 -15.225 4.500 -14.975 ;
        RECT 5.470 -15.185 5.640 -14.895 ;
        RECT 6.440 -15.060 6.610 -14.215 ;
        RECT 7.060 -14.385 7.280 -13.515 ;
        RECT 7.505 -13.635 8.200 -13.445 ;
        RECT 6.780 -14.765 7.280 -14.385 ;
        RECT 7.450 -14.435 7.860 -13.815 ;
        RECT 8.030 -14.605 8.200 -13.635 ;
        RECT 7.505 -14.775 8.200 -14.605 ;
        RECT 6.440 -15.230 7.270 -15.060 ;
        RECT 7.505 -15.275 7.675 -14.775 ;
        RECT 8.390 -15.275 8.615 -13.155 ;
        RECT 9.285 -13.445 9.455 -13.155 ;
        RECT 8.790 -13.615 9.455 -13.445 ;
        RECT 8.790 -14.605 9.020 -13.615 ;
        RECT 12.085 -13.640 12.340 -13.065 ;
        RECT 13.055 -13.445 13.225 -13.065 ;
        RECT 12.510 -13.615 13.225 -13.445 ;
        RECT 9.190 -13.800 9.540 -13.785 ;
        RECT 9.190 -14.150 11.100 -13.800 ;
        RECT 9.190 -14.435 9.540 -14.150 ;
        RECT 12.085 -14.370 12.255 -13.640 ;
        RECT 12.510 -13.805 12.680 -13.615 ;
        RECT 12.425 -14.135 12.680 -13.805 ;
        RECT 12.510 -14.345 12.680 -14.135 ;
        RECT 8.790 -14.775 9.455 -14.605 ;
        RECT 9.285 -15.275 9.455 -14.775 ;
        RECT 12.085 -15.275 12.340 -14.370 ;
        RECT 12.510 -14.515 13.225 -14.345 ;
        RECT 13.055 -15.275 13.225 -14.515 ;
      LAYER met1 ;
        RECT 0.480 -3.220 0.770 -3.175 ;
        RECT 2.340 -3.220 2.630 -3.175 ;
        RECT 5.120 -3.220 5.410 -3.175 ;
        RECT 0.480 -3.360 5.410 -3.220 ;
        RECT 0.480 -3.405 0.770 -3.360 ;
        RECT 2.340 -3.405 2.630 -3.360 ;
        RECT 5.120 -3.405 5.410 -3.360 ;
        RECT 12.450 -3.400 14.750 -3.050 ;
        RECT -1.050 -4.050 2.100 -3.650 ;
        RECT 5.120 -3.900 5.410 -3.855 ;
        RECT 2.875 -4.040 5.410 -3.900 ;
        RECT -2.350 -9.000 -1.900 -8.950 ;
        RECT -2.750 -9.350 -1.900 -9.000 ;
        RECT -2.350 -9.400 -1.900 -9.350 ;
        RECT -1.050 -10.900 -0.700 -4.050 ;
        RECT 2.875 -4.195 3.090 -4.040 ;
        RECT 5.120 -4.085 5.410 -4.040 ;
        RECT 0.940 -4.240 1.230 -4.195 ;
        RECT 2.800 -4.240 3.090 -4.195 ;
        RECT 3.720 -4.200 4.010 -4.195 ;
        RECT 0.940 -4.380 3.090 -4.240 ;
        RECT 0.940 -4.425 1.230 -4.380 ;
        RECT 2.800 -4.425 3.090 -4.380 ;
        RECT 3.650 -4.240 4.150 -4.200 ;
        RECT 6.980 -4.240 7.270 -4.195 ;
        RECT 3.650 -4.380 7.270 -4.240 ;
        RECT 3.650 -4.650 4.150 -4.380 ;
        RECT 6.980 -4.425 7.270 -4.380 ;
        RECT 10.400 -6.650 10.750 -3.800 ;
        RECT 3.050 -7.000 10.750 -6.650 ;
        RECT 3.050 -8.650 3.400 -7.000 ;
        RECT 3.050 -9.000 5.950 -8.650 ;
        RECT 5.000 -9.850 5.350 -9.500 ;
        RECT 5.600 -9.550 5.950 -9.000 ;
        RECT 5.500 -9.800 6.050 -9.550 ;
        RECT -3.700 -11.200 -0.700 -10.900 ;
        RECT 3.050 -10.200 5.350 -9.850 ;
        RECT -3.700 -13.350 -3.350 -11.200 ;
        RECT 3.050 -11.900 3.400 -10.200 ;
        RECT 14.400 -11.700 14.750 -3.400 ;
        RECT -0.700 -12.250 3.400 -11.900 ;
        RECT 10.050 -12.050 14.750 -11.700 ;
        RECT -0.700 -13.300 -0.350 -12.250 ;
        RECT -3.700 -13.700 -1.650 -13.350 ;
        RECT -0.700 -13.700 0.750 -13.300 ;
        RECT 2.290 -13.590 2.580 -13.545 ;
        RECT 5.550 -13.590 6.050 -13.250 ;
        RECT 2.290 -13.730 6.050 -13.590 ;
        RECT 2.290 -13.775 2.580 -13.730 ;
        RECT 5.550 -13.750 6.050 -13.730 ;
        RECT 6.470 -13.590 6.760 -13.545 ;
        RECT 8.330 -13.590 8.620 -13.545 ;
        RECT 6.470 -13.730 8.620 -13.590 ;
        RECT 5.550 -13.775 5.840 -13.750 ;
        RECT 6.470 -13.775 6.760 -13.730 ;
        RECT 8.330 -13.775 8.620 -13.730 ;
        RECT 4.150 -13.930 4.440 -13.885 ;
        RECT 6.470 -13.930 6.685 -13.775 ;
        RECT 4.150 -14.070 6.685 -13.930 ;
        RECT 4.150 -14.115 4.440 -14.070 ;
        RECT 7.450 -14.100 7.850 -13.900 ;
        RECT 10.050 -14.100 10.400 -12.050 ;
        RECT 7.450 -14.400 10.400 -14.100 ;
        RECT 10.750 -14.150 12.400 -13.800 ;
        RECT 7.450 -14.450 8.650 -14.400 ;
        RECT 9.250 -14.450 10.400 -14.400 ;
        RECT 4.150 -14.610 4.440 -14.565 ;
        RECT 6.930 -14.610 7.220 -14.565 ;
        RECT 8.790 -14.610 9.080 -14.565 ;
        RECT 4.150 -14.750 9.080 -14.610 ;
        RECT 4.150 -14.795 4.440 -14.750 ;
        RECT 6.930 -14.795 7.220 -14.750 ;
        RECT 8.790 -14.795 9.080 -14.750 ;
        RECT 12.050 -14.950 12.400 -14.150 ;
      LAYER met2 ;
        RECT 3.650 -4.750 4.150 -4.200 ;
        RECT 3.650 -5.900 4.000 -4.750 ;
        RECT 0.500 -6.250 4.000 -5.900 ;
        RECT -2.350 -9.000 -1.900 -8.950 ;
        RECT 0.500 -9.000 0.850 -6.250 ;
        RECT -2.350 -9.350 0.850 -9.000 ;
        RECT -2.350 -9.400 -1.900 -9.350 ;
        RECT 0.500 -11.300 0.850 -9.350 ;
        RECT 0.500 -11.650 5.900 -11.300 ;
        RECT 5.550 -13.250 5.900 -11.650 ;
        RECT 5.550 -13.750 6.050 -13.250 ;
  END
END count
MACRO dco
  CLASS BLOCK ;
  FOREIGN dco ;
  ORIGIN 3.600 21.400 ;
  SIZE 63.300 BY 52.200 ;
  PIN VCCD
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.917700 ;
    PORT
      LAYER nwell ;
        RECT 15.400 17.500 18.930 19.100 ;
        RECT 16.250 17.495 18.930 17.500 ;
        RECT 33.850 4.500 36.700 6.100 ;
        RECT 33.850 4.495 36.070 4.500 ;
        RECT 39.550 3.400 41.700 3.450 ;
        RECT 39.550 1.800 53.940 3.400 ;
        RECT 41.600 1.795 53.940 1.800 ;
        RECT 44.200 1.750 46.300 1.795 ;
        RECT 38.550 -2.400 56.300 -0.800 ;
        RECT 39.400 -2.405 56.300 -2.400 ;
        RECT 42.500 -2.450 44.850 -2.405 ;
        RECT 54.800 -2.450 56.300 -2.405 ;
        RECT 6.545 -9.700 8.150 -7.550 ;
        RECT 6.500 -10.850 8.150 -9.700 ;
        RECT 39.550 -8.300 41.700 -8.250 ;
        RECT 39.550 -9.900 53.940 -8.300 ;
        RECT 41.600 -9.905 53.940 -9.900 ;
        RECT 44.200 -9.950 46.300 -9.905 ;
        RECT 6.545 -12.610 8.150 -10.850 ;
        RECT 38.550 -14.100 56.300 -12.500 ;
        RECT 39.400 -14.105 56.300 -14.100 ;
        RECT 42.500 -14.150 44.850 -14.105 ;
        RECT 54.800 -14.150 56.300 -14.105 ;
      LAYER li1 ;
        RECT 16.440 18.825 18.740 18.995 ;
        RECT 15.800 17.980 16.100 18.480 ;
        RECT 16.955 18.425 17.890 18.825 ;
        RECT 18.415 17.500 18.655 18.145 ;
        RECT 18.415 17.200 18.800 17.500 ;
        RECT 18.415 17.165 18.655 17.200 ;
        RECT 39.750 6.450 42.300 6.950 ;
        RECT 34.040 5.825 35.880 5.995 ;
        RECT 34.600 5.065 34.930 5.825 ;
        RECT 35.530 4.675 35.790 5.825 ;
        RECT 36.150 4.750 36.450 5.250 ;
        RECT 39.750 2.400 40.250 6.450 ;
        RECT 41.800 3.295 42.300 6.450 ;
        RECT 53.700 3.295 55.050 3.450 ;
        RECT 41.790 3.125 44.090 3.295 ;
        RECT 46.390 3.125 55.050 3.295 ;
        RECT 41.920 1.985 42.185 3.125 ;
        RECT 42.855 2.325 43.025 3.125 ;
        RECT 43.695 2.665 43.905 3.125 ;
        RECT 46.905 2.625 47.235 3.125 ;
        RECT 47.830 2.665 48.095 3.125 ;
        RECT 50.000 2.325 50.170 3.125 ;
        RECT 51.880 2.625 52.195 3.125 ;
        RECT 52.935 2.115 53.105 3.125 ;
        RECT 53.700 3.100 55.050 3.125 ;
        RECT 54.650 -0.650 55.050 3.100 ;
        RECT 42.350 -0.905 44.000 -0.750 ;
        RECT 39.590 -1.075 44.000 -0.905 ;
        RECT 44.990 -1.075 54.650 -0.905 ;
        RECT 38.850 -1.850 39.250 -1.350 ;
        RECT 40.185 -1.875 40.425 -1.075 ;
        RECT 40.945 -1.875 41.275 -1.075 ;
        RECT 41.785 -2.225 42.115 -1.075 ;
        RECT 42.350 -1.200 44.000 -1.075 ;
        RECT 45.505 -1.575 45.835 -1.075 ;
        RECT 46.430 -1.535 46.695 -1.075 ;
        RECT 48.600 -1.875 48.770 -1.075 ;
        RECT 50.480 -1.575 50.795 -1.075 ;
        RECT 51.540 -2.085 51.710 -1.075 ;
        RECT 52.380 -1.990 52.555 -1.075 ;
        RECT 53.415 -2.215 53.630 -1.075 ;
        RECT 54.305 -2.215 54.555 -1.075 ;
        RECT 55.000 -2.200 55.500 -1.800 ;
        RECT 7.875 -8.300 8.045 -7.740 ;
        RECT 7.115 -8.630 8.045 -8.300 ;
        RECT 53.700 -8.405 55.050 -8.250 ;
        RECT 41.790 -8.575 44.090 -8.405 ;
        RECT 46.390 -8.575 55.050 -8.405 ;
        RECT 7.875 -9.230 8.045 -8.630 ;
        RECT 6.725 -9.490 8.045 -9.230 ;
        RECT 39.850 -9.300 40.250 -8.800 ;
        RECT 7.875 -9.580 8.045 -9.490 ;
        RECT 41.920 -9.715 42.185 -8.575 ;
        RECT 42.855 -9.375 43.025 -8.575 ;
        RECT 43.695 -9.035 43.905 -8.575 ;
        RECT 46.905 -9.075 47.235 -8.575 ;
        RECT 47.830 -9.035 48.095 -8.575 ;
        RECT 50.000 -9.375 50.170 -8.575 ;
        RECT 51.880 -9.075 52.195 -8.575 ;
        RECT 52.935 -9.585 53.105 -8.575 ;
        RECT 53.700 -8.600 55.050 -8.575 ;
        RECT 6.900 -10.200 7.400 -9.800 ;
        RECT 7.875 -11.165 8.045 -11.040 ;
        RECT 6.735 -11.395 8.045 -11.165 ;
        RECT 7.875 -12.065 8.045 -11.395 ;
        RECT 6.735 -12.275 8.045 -12.065 ;
        RECT 7.875 -12.420 8.045 -12.275 ;
        RECT 54.650 -12.350 55.050 -8.600 ;
        RECT 42.350 -12.605 44.000 -12.450 ;
        RECT 39.590 -12.775 44.000 -12.605 ;
        RECT 44.990 -12.775 54.650 -12.605 ;
        RECT 38.850 -13.550 39.250 -13.050 ;
        RECT 40.185 -13.575 40.425 -12.775 ;
        RECT 40.945 -13.575 41.275 -12.775 ;
        RECT 41.785 -13.925 42.115 -12.775 ;
        RECT 42.350 -12.900 44.000 -12.775 ;
        RECT 45.505 -13.275 45.835 -12.775 ;
        RECT 46.430 -13.235 46.695 -12.775 ;
        RECT 48.600 -13.575 48.770 -12.775 ;
        RECT 50.480 -13.275 50.795 -12.775 ;
        RECT 51.540 -13.785 51.710 -12.775 ;
        RECT 52.380 -13.690 52.555 -12.775 ;
        RECT 53.415 -13.915 53.630 -12.775 ;
        RECT 54.305 -13.915 54.555 -12.775 ;
        RECT 55.000 -13.900 55.500 -13.500 ;
      LAYER met1 ;
        RECT 15.800 18.700 18.740 19.150 ;
        RECT 15.800 17.980 16.100 18.700 ;
        RECT 16.440 18.670 18.740 18.700 ;
        RECT 19.600 17.500 20.050 19.150 ;
        RECT 18.400 17.150 20.050 17.500 ;
        RECT 35.900 6.150 36.450 6.950 ;
        RECT 39.750 6.450 42.300 6.950 ;
        RECT 34.040 5.700 36.450 6.150 ;
        RECT 34.040 5.670 35.880 5.700 ;
        RECT 36.150 4.750 36.450 5.700 ;
        RECT 41.790 2.970 53.750 3.450 ;
        RECT 44.050 2.950 46.500 2.970 ;
        RECT 38.000 2.400 40.250 2.900 ;
        RECT 38.000 -1.350 38.500 2.400 ;
        RECT 54.650 -0.750 55.050 -0.250 ;
        RECT 39.590 -1.230 42.350 -0.750 ;
        RECT 43.500 -1.200 55.050 -0.750 ;
        RECT 44.990 -1.230 55.050 -1.200 ;
        RECT 54.650 -1.250 55.050 -1.230 ;
        RECT 38.000 -1.850 39.250 -1.350 ;
        RECT 55.000 -2.200 55.500 -1.800 ;
        RECT 7.700 -7.750 8.200 -6.700 ;
        RECT 7.720 -9.550 8.200 -7.750 ;
        RECT 41.790 -8.730 53.750 -8.250 ;
        RECT 44.050 -8.750 46.500 -8.730 ;
        RECT 32.650 -9.300 40.250 -8.800 ;
        RECT 7.700 -9.800 8.200 -9.550 ;
        RECT 6.900 -10.200 8.200 -9.800 ;
        RECT 7.700 -11.050 8.200 -10.200 ;
        RECT 7.720 -12.420 8.200 -11.050 ;
        RECT 38.000 -12.450 38.500 -9.300 ;
        RECT 54.650 -12.450 55.050 -11.950 ;
        RECT 38.000 -12.900 42.350 -12.450 ;
        RECT 43.500 -12.900 55.050 -12.450 ;
        RECT 38.000 -13.050 38.500 -12.900 ;
        RECT 39.590 -12.930 42.350 -12.900 ;
        RECT 44.990 -12.930 55.050 -12.900 ;
        RECT 54.650 -12.950 55.050 -12.930 ;
        RECT 38.000 -13.550 39.250 -13.050 ;
        RECT 55.000 -13.900 55.500 -13.500 ;
      LAYER met2 ;
        RECT -3.600 19.150 -2.650 30.400 ;
        RECT -3.600 18.700 20.050 19.150 ;
        RECT -3.600 6.950 -2.650 18.700 ;
        RECT -3.600 6.500 42.300 6.950 ;
        RECT -3.600 0.725 -2.650 6.500 ;
        RECT 7.700 -7.200 8.200 6.500 ;
        RECT 32.650 -9.300 33.150 6.500 ;
        RECT 39.750 6.450 42.300 6.500 ;
    END
  END VCCD
  PIN VCCA
    ANTENNADIFFAREA 2.560000 ;
    PORT
      LAYER nwell ;
        RECT 11.400 -0.700 13.800 1.900 ;
        RECT 15.150 -0.700 19.350 1.900 ;
      LAYER li1 ;
        RECT 10.800 3.000 18.250 3.400 ;
        RECT 11.600 1.000 12.000 3.000 ;
        RECT 12.300 -0.300 12.700 3.000 ;
        RECT 15.350 1.050 15.750 3.000 ;
        RECT 16.050 -0.300 16.450 1.500 ;
        RECT 17.850 -0.300 18.250 3.000 ;
      LAYER met1 ;
        RECT 11.600 1.000 12.000 1.500 ;
        RECT 15.350 1.050 15.750 1.550 ;
        RECT 16.050 1.350 16.450 1.500 ;
        RECT 17.850 1.350 18.250 1.500 ;
        RECT 16.050 0.850 18.250 1.350 ;
        RECT 16.050 0.700 16.450 0.850 ;
        RECT 17.850 0.700 18.250 0.850 ;
    END
  END VCCA
  PIN Dctrl
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 6.225 -8.180 6.595 -7.825 ;
      LAYER met1 ;
        RECT 6.200 -8.200 6.600 -6.700 ;
    END
  END Dctrl
  PIN ENB
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 16.525 17.185 16.985 17.915 ;
      LAYER met1 ;
        RECT 16.500 17.450 17.000 17.700 ;
        RECT 14.450 17.150 17.000 17.450 ;
    END
  END ENB
  PIN Vbs_12
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 12.900 1.900 13.200 2.400 ;
        RECT 27.450 1.850 27.950 2.350 ;
      LAYER met1 ;
        RECT 12.700 4.350 13.200 4.800 ;
        RECT 12.700 3.850 27.950 4.350 ;
        RECT 12.700 1.900 13.200 3.850 ;
        RECT 27.450 1.850 27.950 3.850 ;
    END
  END Vbs_12
  PIN Vbs_34
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER li1 ;
        RECT 16.650 1.900 17.650 2.400 ;
        RECT 21.950 1.900 24.250 2.400 ;
      LAYER met1 ;
        RECT 19.800 2.400 20.300 2.950 ;
        RECT 16.450 1.900 24.250 2.400 ;
    END
  END Vbs_34
  PIN pha_DCO
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 51.880 -13.835 52.210 -12.990 ;
        RECT 51.880 -13.915 52.290 -13.835 ;
        RECT 52.055 -13.965 52.290 -13.915 ;
        RECT 52.100 -14.545 52.290 -13.965 ;
        RECT 52.045 -14.585 52.290 -14.545 ;
        RECT 51.890 -14.670 52.290 -14.585 ;
        RECT 51.890 -15.105 52.220 -14.670 ;
      LAYER met1 ;
        RECT 55.400 -13.100 55.900 -11.950 ;
        RECT 51.850 -13.350 55.900 -13.100 ;
        RECT 51.850 -14.150 52.300 -13.350 ;
        RECT 51.850 -14.900 52.350 -14.150 ;
      LAYER met2 ;
        RECT 55.400 -12.450 59.450 -11.950 ;
    END
  END pha_DCO
  PIN GND
    ANTENNADIFFAREA 42.328999 ;
    PORT
      LAYER pwell ;
        RECT 8.400 21.800 51.600 24.600 ;
        RECT 16.930 16.975 18.735 17.205 ;
        RECT 16.445 16.970 18.735 16.975 ;
        RECT 15.780 16.295 18.735 16.970 ;
        RECT 15.780 16.290 16.450 16.295 ;
        RECT 16.590 16.105 16.760 16.295 ;
        RECT 22.850 13.600 51.650 16.400 ;
        RECT 34.530 4.200 35.875 4.205 ;
        RECT 34.530 3.975 36.700 4.200 ;
        RECT 34.045 3.300 36.700 3.975 ;
        RECT 34.045 3.295 35.875 3.300 ;
        RECT 34.185 3.105 34.355 3.295 ;
        RECT 39.550 1.505 41.900 1.550 ;
        RECT 39.550 1.300 44.035 1.505 ;
        RECT 39.550 1.275 46.450 1.300 ;
        RECT 49.910 1.275 50.820 1.495 ;
        RECT 52.355 1.275 53.705 1.505 ;
        RECT 39.550 0.595 53.705 1.275 ;
        RECT 39.550 0.550 41.900 0.595 ;
        RECT 41.935 0.405 42.105 0.595 ;
        RECT 44.000 0.550 46.450 0.595 ;
        RECT 46.535 0.405 46.705 0.595 ;
        RECT 39.595 -2.700 42.205 -2.695 ;
        RECT 38.550 -2.900 42.205 -2.700 ;
        RECT 38.550 -2.925 45.050 -2.900 ;
        RECT 48.510 -2.925 49.420 -2.705 ;
        RECT 50.960 -2.925 54.645 -2.695 ;
        RECT 38.550 -3.605 54.645 -2.925 ;
        RECT 38.550 -3.950 39.650 -3.605 ;
        RECT 39.740 -3.795 39.910 -3.605 ;
        RECT 42.200 -3.650 45.050 -3.605 ;
        RECT 45.135 -3.795 45.305 -3.605 ;
        RECT 5.345 -7.885 6.025 -7.745 ;
        RECT 5.155 -8.055 6.025 -7.885 ;
        RECT 5.345 -8.230 6.025 -8.055 ;
        RECT 16.550 -8.100 19.850 -5.300 ;
        RECT 21.100 -8.100 24.400 -5.300 ;
        RECT 5.345 -9.575 6.255 -8.230 ;
        RECT 5.350 -11.055 6.250 -9.575 ;
        RECT 39.550 -10.195 41.900 -10.150 ;
        RECT 39.550 -10.400 44.035 -10.195 ;
        RECT 39.550 -10.425 46.450 -10.400 ;
        RECT 49.910 -10.425 50.820 -10.205 ;
        RECT 52.355 -10.425 53.705 -10.195 ;
        RECT 5.345 -11.185 6.255 -11.055 ;
        RECT 39.550 -11.105 53.705 -10.425 ;
        RECT 39.550 -11.150 41.900 -11.105 ;
        RECT 5.155 -11.355 6.255 -11.185 ;
        RECT 41.935 -11.295 42.105 -11.105 ;
        RECT 44.000 -11.150 46.450 -11.105 ;
        RECT 46.535 -11.295 46.705 -11.105 ;
        RECT 5.345 -12.405 6.255 -11.355 ;
        RECT 14.000 -16.100 28.380 -14.090 ;
        RECT 39.595 -14.400 42.205 -14.395 ;
        RECT 38.550 -14.600 42.205 -14.400 ;
        RECT 38.550 -14.625 45.050 -14.600 ;
        RECT 48.510 -14.625 49.420 -14.405 ;
        RECT 50.960 -14.625 54.645 -14.395 ;
        RECT 38.550 -15.305 54.645 -14.625 ;
        RECT 38.550 -15.650 39.650 -15.305 ;
        RECT 39.740 -15.495 39.910 -15.305 ;
        RECT 42.200 -15.350 45.050 -15.305 ;
        RECT 45.135 -15.495 45.305 -15.305 ;
      LAYER li1 ;
        RECT 8.600 22.150 9.000 22.650 ;
        RECT 9.300 21.300 9.700 24.200 ;
        RECT 12.100 21.300 12.500 24.200 ;
        RECT 12.900 22.150 13.300 22.650 ;
        RECT 13.600 21.300 14.000 24.200 ;
        RECT 15.800 22.150 16.200 22.650 ;
        RECT 16.500 21.300 16.900 24.200 ;
        RECT 18.700 22.150 19.100 22.650 ;
        RECT 19.400 21.300 19.800 24.200 ;
        RECT 22.200 21.300 22.600 24.200 ;
        RECT 23.000 22.150 23.400 22.650 ;
        RECT 23.700 21.300 24.100 24.200 ;
        RECT 26.500 21.300 26.900 24.200 ;
        RECT 27.300 22.150 27.700 22.650 ;
        RECT 28.000 21.300 28.400 24.200 ;
        RECT 30.200 22.150 30.600 22.650 ;
        RECT 30.900 21.300 31.300 24.200 ;
        RECT 33.100 22.150 33.500 22.650 ;
        RECT 33.800 21.300 34.200 24.200 ;
        RECT 36.600 21.300 37.000 24.200 ;
        RECT 37.400 22.150 37.800 22.650 ;
        RECT 38.100 21.300 38.500 24.200 ;
        RECT 40.900 21.300 41.300 24.200 ;
        RECT 41.700 22.150 42.100 22.650 ;
        RECT 42.400 21.300 42.800 24.200 ;
        RECT 44.600 22.150 45.000 22.650 ;
        RECT 45.300 21.300 45.700 24.200 ;
        RECT 47.500 22.150 47.900 22.650 ;
        RECT 48.200 21.300 48.600 24.200 ;
        RECT 51.000 21.300 51.400 24.200 ;
        RECT 9.300 20.900 51.400 21.300 ;
        RECT 23.050 17.300 23.450 20.900 ;
        RECT 50.350 17.300 50.750 20.900 ;
        RECT 22.000 16.900 50.750 17.300 ;
        RECT 15.850 15.850 16.200 16.900 ;
        RECT 16.955 16.275 17.890 16.675 ;
        RECT 16.440 16.105 18.740 16.275 ;
        RECT 16.450 15.850 16.800 16.105 ;
        RECT 15.850 15.500 16.800 15.850 ;
        RECT 15.850 13.650 16.350 15.500 ;
        RECT 22.000 13.650 22.400 16.900 ;
        RECT 23.050 14.000 23.450 16.900 ;
        RECT 25.850 14.000 26.250 16.900 ;
        RECT 26.550 15.550 26.950 16.050 ;
        RECT 28.750 14.000 29.150 16.900 ;
        RECT 29.450 15.550 29.850 16.050 ;
        RECT 31.650 14.000 32.050 16.900 ;
        RECT 32.350 15.550 32.750 16.050 ;
        RECT 33.150 14.000 33.550 16.900 ;
        RECT 35.950 14.000 36.350 16.900 ;
        RECT 36.650 15.550 37.050 16.050 ;
        RECT 37.450 14.000 37.850 16.900 ;
        RECT 40.250 14.000 40.650 16.900 ;
        RECT 40.950 15.550 41.350 16.050 ;
        RECT 43.150 14.000 43.550 16.900 ;
        RECT 43.850 15.550 44.250 16.050 ;
        RECT 46.050 14.000 46.450 16.900 ;
        RECT 46.750 15.550 47.150 16.050 ;
        RECT 47.550 14.000 47.950 16.900 ;
        RECT 50.350 14.000 50.750 16.900 ;
        RECT 51.050 15.550 51.450 16.050 ;
        RECT 15.850 13.250 22.400 13.650 ;
        RECT 15.850 4.700 16.350 13.250 ;
        RECT 34.600 3.275 34.930 3.655 ;
        RECT 35.530 3.275 35.790 4.115 ;
        RECT 34.040 3.105 35.880 3.275 ;
        RECT 35.450 2.450 35.850 3.105 ;
        RECT 36.150 2.450 36.450 4.000 ;
        RECT 35.450 2.150 36.450 2.450 ;
        RECT 35.450 1.250 35.850 2.150 ;
        RECT 35.450 0.750 40.250 1.250 ;
        RECT 35.450 0.550 35.950 0.750 ;
        RECT 41.920 0.600 42.185 1.035 ;
        RECT 41.920 0.575 42.200 0.600 ;
        RECT 42.855 0.575 43.025 1.035 ;
        RECT 43.695 0.575 43.945 1.040 ;
        RECT 46.905 0.575 47.235 0.955 ;
        RECT 47.845 0.575 48.095 1.035 ;
        RECT 49.790 0.575 50.160 1.075 ;
        RECT 51.975 0.575 52.185 1.105 ;
        RECT 52.945 0.575 53.115 1.185 ;
        RECT 41.790 0.550 44.090 0.575 ;
        RECT 35.450 0.405 44.090 0.550 ;
        RECT 46.390 0.405 53.750 0.575 ;
        RECT 35.450 0.150 42.200 0.405 ;
        RECT 16.750 -6.150 17.150 -5.650 ;
        RECT 5.155 -8.300 5.325 -7.740 ;
        RECT 23.800 -7.750 24.200 -7.250 ;
        RECT 5.155 -8.630 5.705 -8.300 ;
        RECT 5.155 -9.230 5.325 -8.630 ;
        RECT 5.155 -9.490 6.165 -9.230 ;
        RECT 5.155 -9.580 5.325 -9.490 ;
        RECT 5.500 -10.300 6.000 -9.900 ;
        RECT 35.450 -10.450 35.950 0.150 ;
        RECT 38.850 -3.650 39.250 -3.150 ;
        RECT 40.115 -3.625 40.355 -3.145 ;
        RECT 40.945 -3.625 41.275 -3.145 ;
        RECT 41.785 -3.625 42.115 -2.825 ;
        RECT 42.350 -3.625 45.000 -3.450 ;
        RECT 45.505 -3.625 45.835 -3.245 ;
        RECT 46.445 -3.625 46.695 -3.165 ;
        RECT 48.390 -3.625 48.760 -3.125 ;
        RECT 50.575 -3.625 50.785 -3.095 ;
        RECT 51.550 -3.625 51.720 -3.015 ;
        RECT 52.390 -3.625 52.560 -3.110 ;
        RECT 53.380 -3.625 53.710 -2.885 ;
        RECT 54.305 -3.625 54.555 -2.805 ;
        RECT 39.590 -3.795 54.650 -3.625 ;
        RECT 42.350 -3.950 45.000 -3.795 ;
        RECT 35.450 -10.950 40.250 -10.450 ;
        RECT 5.155 -11.165 5.325 -11.040 ;
        RECT 35.450 -11.150 35.950 -10.950 ;
        RECT 41.920 -11.100 42.185 -10.665 ;
        RECT 41.920 -11.125 42.250 -11.100 ;
        RECT 42.855 -11.125 43.025 -10.665 ;
        RECT 43.695 -11.125 43.945 -10.660 ;
        RECT 46.905 -11.125 47.235 -10.745 ;
        RECT 47.845 -11.125 48.095 -10.665 ;
        RECT 49.790 -11.125 50.160 -10.625 ;
        RECT 51.975 -11.125 52.185 -10.595 ;
        RECT 52.945 -11.125 53.115 -10.515 ;
        RECT 41.790 -11.150 44.090 -11.125 ;
        RECT 5.155 -11.395 6.145 -11.165 ;
        RECT 35.450 -11.295 44.090 -11.150 ;
        RECT 46.390 -11.295 53.750 -11.125 ;
        RECT 5.155 -12.065 5.325 -11.395 ;
        RECT 35.450 -11.500 42.250 -11.295 ;
        RECT 5.155 -12.275 6.145 -12.065 ;
        RECT 5.155 -12.420 5.325 -12.275 ;
        RECT 12.300 -13.600 17.150 -13.200 ;
        RECT 14.180 -14.440 28.200 -14.270 ;
        RECT 14.180 -15.600 14.350 -14.440 ;
        RECT 27.450 -14.920 27.750 -14.900 ;
        RECT 25.390 -15.270 27.750 -14.920 ;
        RECT 13.750 -15.750 14.750 -15.600 ;
        RECT 27.450 -15.750 27.750 -15.270 ;
        RECT 28.030 -15.750 28.200 -14.440 ;
        RECT 13.750 -15.920 28.200 -15.750 ;
        RECT 13.750 -20.400 14.750 -15.920 ;
        RECT 35.450 -20.400 35.950 -11.500 ;
        RECT 38.850 -15.350 39.250 -14.850 ;
        RECT 40.115 -15.325 40.355 -14.845 ;
        RECT 40.945 -15.325 41.275 -14.845 ;
        RECT 41.785 -15.325 42.115 -14.525 ;
        RECT 42.350 -15.325 45.000 -15.150 ;
        RECT 45.505 -15.325 45.835 -14.945 ;
        RECT 46.445 -15.325 46.695 -14.865 ;
        RECT 48.390 -15.325 48.760 -14.825 ;
        RECT 50.575 -15.325 50.785 -14.795 ;
        RECT 51.550 -15.325 51.720 -14.715 ;
        RECT 52.390 -15.325 52.560 -14.810 ;
        RECT 53.380 -15.325 53.710 -14.585 ;
        RECT 54.305 -15.325 54.555 -14.505 ;
        RECT 39.590 -15.495 54.650 -15.325 ;
        RECT 42.350 -15.650 45.000 -15.495 ;
        RECT 13.750 -21.400 37.100 -20.400 ;
      LAYER met1 ;
        RECT 8.600 20.400 9.000 22.650 ;
        RECT 12.900 20.400 13.300 22.650 ;
        RECT 15.800 20.400 16.200 22.650 ;
        RECT 18.700 20.400 19.100 22.650 ;
        RECT 23.000 20.400 23.400 22.650 ;
        RECT 27.300 20.400 27.700 22.650 ;
        RECT 30.200 20.400 30.600 22.650 ;
        RECT 33.100 20.400 33.500 22.650 ;
        RECT 37.400 20.400 37.800 22.650 ;
        RECT 41.700 20.400 42.100 22.650 ;
        RECT 44.600 20.400 45.000 22.650 ;
        RECT 47.500 20.400 47.900 22.650 ;
        RECT 8.600 20.000 47.900 20.400 ;
        RECT 26.550 18.200 26.950 20.000 ;
        RECT 47.500 18.200 47.900 20.000 ;
        RECT 26.550 17.800 51.450 18.200 ;
        RECT 15.890 16.380 16.200 16.880 ;
        RECT 16.440 15.950 18.740 16.430 ;
        RECT 26.550 15.550 26.950 17.800 ;
        RECT 29.450 15.550 29.850 17.800 ;
        RECT 32.350 15.550 32.750 17.800 ;
        RECT 36.650 15.550 37.050 17.800 ;
        RECT 40.950 15.550 41.350 17.800 ;
        RECT 43.850 15.550 44.250 17.800 ;
        RECT 46.750 15.550 47.150 17.800 ;
        RECT 51.050 15.550 51.450 17.800 ;
        RECT 15.850 4.700 31.350 5.200 ;
        RECT 30.850 1.250 31.350 4.700 ;
        RECT 36.150 3.500 36.450 4.000 ;
        RECT 34.040 2.950 35.880 3.430 ;
        RECT 30.850 0.750 37.700 1.250 ;
        RECT 39.850 0.750 40.250 1.250 ;
        RECT 37.200 -3.150 37.700 0.750 ;
        RECT 41.790 0.600 44.090 0.730 ;
        RECT 46.390 0.650 53.750 0.730 ;
        RECT 46.390 0.600 57.050 0.650 ;
        RECT 41.790 0.250 57.050 0.600 ;
        RECT 37.200 -3.650 39.250 -3.150 ;
        RECT 39.590 -3.950 42.350 -3.470 ;
        RECT 44.990 -3.500 54.650 -3.470 ;
        RECT 56.600 -3.500 57.050 0.250 ;
        RECT 44.990 -3.950 57.050 -3.500 ;
        RECT 5.000 -9.550 5.480 -7.740 ;
        RECT 5.000 -9.900 5.500 -9.550 ;
        RECT 16.750 -9.650 17.150 -5.650 ;
        RECT 23.800 -9.650 24.200 -7.250 ;
        RECT 5.000 -10.300 6.000 -9.900 ;
        RECT 16.750 -10.050 24.200 -9.650 ;
        RECT 5.000 -11.050 5.500 -10.300 ;
        RECT 5.000 -12.420 5.480 -11.050 ;
        RECT 5.050 -15.600 5.450 -12.420 ;
        RECT 12.300 -15.600 12.700 -13.200 ;
        RECT 16.750 -13.600 17.150 -10.050 ;
        RECT 37.200 -14.850 37.700 -10.450 ;
        RECT 39.850 -10.950 40.250 -10.450 ;
        RECT 41.790 -11.100 44.090 -10.970 ;
        RECT 46.390 -11.050 53.750 -10.970 ;
        RECT 46.390 -11.100 57.050 -11.050 ;
        RECT 41.790 -11.450 57.050 -11.100 ;
        RECT 25.415 -15.220 27.520 -14.970 ;
        RECT 37.200 -15.350 39.250 -14.850 ;
        RECT 5.050 -16.000 14.500 -15.600 ;
        RECT 39.590 -15.650 42.350 -15.170 ;
        RECT 44.990 -15.200 54.650 -15.170 ;
        RECT 56.600 -15.200 57.050 -11.450 ;
        RECT 44.990 -15.650 57.050 -15.200 ;
    END
  END GND
  OBS
      LAYER nwell ;
        RECT 8.400 24.900 51.600 28.700 ;
        RECT 22.850 9.500 51.650 13.300 ;
        RECT 20.650 -0.700 24.850 1.900 ;
        RECT 26.150 -0.750 28.550 1.850 ;
      LAYER pwell ;
        RECT 54.650 -3.650 56.300 -2.700 ;
      LAYER nwell ;
        RECT 11.750 -9.950 15.050 -5.150 ;
        RECT 25.600 -10.000 28.900 -5.200 ;
      LAYER pwell ;
        RECT 54.650 -15.350 56.300 -14.400 ;
      LAYER li1 ;
        RECT 9.300 29.200 53.200 29.600 ;
        RECT 8.600 27.850 9.000 28.350 ;
        RECT 9.300 25.300 9.700 29.200 ;
        RECT 9.950 24.500 10.400 24.950 ;
        RECT 10.700 22.200 11.100 28.300 ;
        RECT 12.100 25.300 12.500 29.200 ;
        RECT 12.900 27.750 13.300 28.250 ;
        RECT 13.600 25.300 14.000 29.200 ;
        RECT 15.000 24.950 15.400 28.300 ;
        RECT 15.800 27.750 16.200 28.250 ;
        RECT 16.500 25.300 16.900 29.200 ;
        RECT 11.350 24.500 11.800 24.950 ;
        RECT 14.250 24.550 14.650 24.950 ;
        RECT 15.000 24.550 17.550 24.950 ;
        RECT 15.000 22.200 15.400 24.550 ;
        RECT 17.900 22.200 18.300 28.300 ;
        RECT 18.700 27.850 19.100 28.350 ;
        RECT 19.400 25.300 19.800 29.200 ;
        RECT 20.050 24.500 20.500 24.950 ;
        RECT 20.800 22.200 21.200 28.300 ;
        RECT 22.200 25.300 22.600 29.200 ;
        RECT 23.000 27.850 23.400 28.350 ;
        RECT 23.700 25.300 24.100 29.200 ;
        RECT 21.450 24.500 21.900 24.950 ;
        RECT 24.350 24.500 24.800 24.950 ;
        RECT 25.100 22.200 25.500 28.300 ;
        RECT 26.500 25.300 26.900 29.200 ;
        RECT 27.300 27.750 27.700 28.250 ;
        RECT 28.000 25.300 28.400 29.200 ;
        RECT 29.400 24.950 29.800 28.300 ;
        RECT 30.200 27.750 30.600 28.250 ;
        RECT 30.900 25.300 31.300 29.200 ;
        RECT 25.750 24.500 26.200 24.950 ;
        RECT 28.650 24.550 29.050 24.950 ;
        RECT 29.400 24.550 31.950 24.950 ;
        RECT 29.400 22.200 29.800 24.550 ;
        RECT 32.300 22.200 32.700 28.300 ;
        RECT 33.100 27.850 33.500 28.350 ;
        RECT 33.800 25.300 34.200 29.200 ;
        RECT 34.450 24.500 34.900 24.950 ;
        RECT 35.200 22.200 35.600 28.300 ;
        RECT 36.600 25.300 37.000 29.200 ;
        RECT 37.400 27.850 37.800 28.350 ;
        RECT 38.100 25.300 38.500 29.200 ;
        RECT 35.850 24.500 36.300 24.950 ;
        RECT 38.750 24.500 39.200 24.950 ;
        RECT 39.500 22.200 39.900 28.300 ;
        RECT 40.900 25.300 41.300 29.200 ;
        RECT 41.700 27.750 42.100 28.250 ;
        RECT 42.400 25.300 42.800 29.200 ;
        RECT 43.800 24.950 44.200 28.300 ;
        RECT 44.600 27.750 45.000 28.250 ;
        RECT 45.300 25.300 45.700 29.200 ;
        RECT 40.150 24.500 40.600 24.950 ;
        RECT 43.050 24.550 43.450 24.950 ;
        RECT 43.800 24.550 46.350 24.950 ;
        RECT 43.800 22.200 44.200 24.550 ;
        RECT 46.700 22.200 47.100 28.300 ;
        RECT 47.500 27.850 47.900 28.350 ;
        RECT 48.200 25.300 48.600 29.200 ;
        RECT 48.850 24.500 49.300 24.950 ;
        RECT 49.600 22.200 50.000 28.300 ;
        RECT 51.000 25.300 51.400 29.200 ;
        RECT 50.250 24.500 50.700 24.950 ;
        RECT 16.525 18.255 16.785 18.655 ;
        RECT 18.060 18.650 18.655 18.655 ;
        RECT 18.060 18.350 20.950 18.650 ;
        RECT 18.060 18.315 18.655 18.350 ;
        RECT 16.525 18.085 17.890 18.255 ;
        RECT 17.155 17.015 17.890 18.085 ;
        RECT 16.525 16.845 17.890 17.015 ;
        RECT 18.060 16.995 18.235 18.315 ;
        RECT 16.525 16.445 16.785 16.845 ;
        RECT 18.060 16.445 18.655 16.995 ;
        RECT 20.650 15.200 20.950 18.350 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 23.750 13.250 24.200 13.700 ;
        RECT 23.050 9.000 23.450 12.900 ;
        RECT 24.450 9.900 24.850 16.000 ;
        RECT 25.150 13.250 25.600 13.700 ;
        RECT 25.850 9.000 26.250 12.900 ;
        RECT 26.550 9.850 26.950 10.350 ;
        RECT 27.350 9.900 27.750 16.000 ;
        RECT 30.250 13.650 30.650 16.000 ;
        RECT 28.100 13.250 30.650 13.650 ;
        RECT 31.000 13.250 31.400 13.650 ;
        RECT 33.850 13.250 34.300 13.700 ;
        RECT 28.750 9.000 29.150 12.900 ;
        RECT 29.450 9.950 29.850 10.450 ;
        RECT 30.250 9.900 30.650 13.250 ;
        RECT 31.650 9.000 32.050 12.900 ;
        RECT 32.350 9.950 32.750 10.450 ;
        RECT 33.150 9.000 33.550 12.900 ;
        RECT 34.550 9.900 34.950 16.000 ;
        RECT 35.250 13.250 35.700 13.700 ;
        RECT 38.150 13.250 38.600 13.700 ;
        RECT 35.950 9.000 36.350 12.900 ;
        RECT 36.650 9.850 37.050 10.350 ;
        RECT 37.450 9.000 37.850 12.900 ;
        RECT 38.850 9.900 39.250 16.000 ;
        RECT 39.550 13.250 40.000 13.700 ;
        RECT 40.250 9.000 40.650 12.900 ;
        RECT 40.950 9.850 41.350 10.350 ;
        RECT 41.750 9.900 42.150 16.000 ;
        RECT 44.650 13.650 45.050 16.000 ;
        RECT 42.500 13.250 45.050 13.650 ;
        RECT 45.400 13.250 45.800 13.650 ;
        RECT 48.250 13.250 48.700 13.700 ;
        RECT 43.150 9.000 43.550 12.900 ;
        RECT 43.850 9.950 44.250 10.450 ;
        RECT 44.650 9.900 45.050 13.250 ;
        RECT 46.050 9.000 46.450 12.900 ;
        RECT 46.750 9.950 47.150 10.450 ;
        RECT 47.550 9.000 47.950 12.900 ;
        RECT 48.950 9.900 49.350 16.000 ;
        RECT 49.650 13.250 50.100 13.700 ;
        RECT 50.350 9.000 50.750 12.900 ;
        RECT 51.050 9.850 51.450 10.350 ;
        RECT 52.800 9.000 53.200 29.200 ;
        RECT 23.050 8.600 53.200 9.000 ;
        RECT 13.200 -0.300 13.600 1.500 ;
        RECT 16.950 -0.300 17.350 1.500 ;
        RECT 18.750 -1.050 19.150 1.500 ;
        RECT 20.850 -1.050 21.250 1.550 ;
        RECT 21.550 -1.050 21.950 1.500 ;
        RECT 18.750 -1.450 21.950 -1.050 ;
        RECT 22.450 -3.000 22.850 1.500 ;
        RECT 23.350 -0.300 23.750 1.500 ;
        RECT 24.250 -0.300 24.650 1.500 ;
        RECT 26.350 1.000 26.750 1.500 ;
        RECT 27.050 -0.350 27.450 1.450 ;
        RECT 27.950 0.150 28.350 1.450 ;
        RECT 29.900 0.150 30.400 7.800 ;
        RECT 34.215 4.895 34.385 5.655 ;
        RECT 34.215 4.725 34.930 4.895 ;
        RECT 35.100 4.750 35.355 5.655 ;
        RECT 34.125 4.175 34.480 4.545 ;
        RECT 34.760 4.515 34.930 4.725 ;
        RECT 34.760 4.185 35.015 4.515 ;
        RECT 34.760 3.995 34.930 4.185 ;
        RECT 35.185 4.020 35.355 4.750 ;
        RECT 34.215 3.825 34.930 3.995 ;
        RECT 34.215 3.445 34.385 3.825 ;
        RECT 35.100 3.445 35.355 4.020 ;
        RECT 42.355 2.155 42.685 2.955 ;
        RECT 43.195 2.175 43.525 2.955 ;
        RECT 46.565 2.455 46.735 2.955 ;
        RECT 46.565 2.285 47.230 2.455 ;
        RECT 43.195 2.155 43.960 2.175 ;
        RECT 42.355 2.100 43.960 2.155 ;
        RECT 46.480 2.100 46.830 2.115 ;
        RECT 42.355 1.985 46.830 2.100 ;
        RECT 41.895 1.565 43.525 1.815 ;
        RECT 43.695 1.700 46.830 1.985 ;
        RECT 43.695 1.395 43.960 1.700 ;
        RECT 46.480 1.465 46.830 1.700 ;
        RECT 42.355 1.215 43.960 1.395 ;
        RECT 47.000 1.295 47.230 2.285 ;
        RECT 42.355 0.745 42.685 1.215 ;
        RECT 43.195 0.745 43.525 1.215 ;
        RECT 45.000 0.800 45.550 1.250 ;
        RECT 46.565 1.125 47.230 1.295 ;
        RECT 46.565 0.835 46.735 1.125 ;
        RECT 47.405 0.835 47.590 2.955 ;
        RECT 48.265 2.530 48.515 2.955 ;
        RECT 48.725 2.680 49.830 2.850 ;
        RECT 48.210 2.400 48.515 2.530 ;
        RECT 47.760 1.205 48.040 2.155 ;
        RECT 48.210 1.295 48.380 2.400 ;
        RECT 48.550 1.615 48.790 2.210 ;
        RECT 48.960 2.145 49.490 2.510 ;
        RECT 48.960 1.445 49.130 2.145 ;
        RECT 49.660 2.065 49.830 2.680 ;
        RECT 50.340 2.625 50.590 2.955 ;
        RECT 50.815 2.655 51.700 2.825 ;
        RECT 49.660 1.975 50.170 2.065 ;
        RECT 48.210 1.165 48.435 1.295 ;
        RECT 48.605 1.225 49.130 1.445 ;
        RECT 49.300 1.805 50.170 1.975 ;
        RECT 48.265 1.025 48.435 1.165 ;
        RECT 49.300 1.025 49.470 1.805 ;
        RECT 50.000 1.735 50.170 1.805 ;
        RECT 49.680 1.555 49.880 1.585 ;
        RECT 50.340 1.555 50.510 2.625 ;
        RECT 50.680 1.735 50.870 2.455 ;
        RECT 49.680 1.255 50.510 1.555 ;
        RECT 51.040 1.525 51.360 2.485 ;
        RECT 48.265 0.855 48.600 1.025 ;
        RECT 48.795 0.855 49.470 1.025 ;
        RECT 50.340 1.025 50.510 1.255 ;
        RECT 50.895 1.195 51.360 1.525 ;
        RECT 51.530 1.815 51.700 2.655 ;
        RECT 52.425 2.395 52.765 2.955 ;
        RECT 51.870 2.020 52.765 2.395 ;
        RECT 52.575 1.815 52.765 2.020 ;
        RECT 53.275 2.065 53.605 2.910 ;
        RECT 53.275 1.985 53.665 2.065 ;
        RECT 53.450 1.935 53.665 1.985 ;
        RECT 51.530 1.485 52.405 1.815 ;
        RECT 52.575 1.485 53.325 1.815 ;
        RECT 51.530 1.025 51.700 1.485 ;
        RECT 52.575 1.315 52.775 1.485 ;
        RECT 53.495 1.355 53.665 1.935 ;
        RECT 53.440 1.315 53.665 1.355 ;
        RECT 50.340 0.855 50.745 1.025 ;
        RECT 50.915 0.855 51.700 1.025 ;
        RECT 27.950 -0.350 30.400 0.150 ;
        RECT 45.175 -0.075 45.425 0.800 ;
        RECT 52.445 0.790 52.775 1.315 ;
        RECT 53.285 1.230 53.665 1.315 ;
        RECT 53.285 0.795 53.615 1.230 ;
        RECT 14.350 -3.500 26.200 -3.000 ;
        RECT 14.350 -4.000 14.850 -3.500 ;
        RECT 11.950 -4.500 14.850 -4.000 ;
        RECT 11.950 -6.000 12.350 -4.500 ;
        RECT 5.495 -8.085 6.045 -7.915 ;
        RECT 5.875 -8.460 6.045 -8.085 ;
        RECT 6.775 -8.085 7.705 -7.915 ;
        RECT 6.775 -8.460 6.945 -8.085 ;
        RECT 5.875 -8.630 6.945 -8.460 ;
        RECT 6.235 -8.715 6.565 -8.630 ;
        RECT 5.495 -8.885 6.070 -8.800 ;
        RECT 6.800 -8.885 7.705 -8.800 ;
        RECT 5.495 -9.055 7.705 -8.885 ;
        RECT 6.350 -10.400 6.550 -9.055 ;
        RECT 12.650 -9.550 13.050 -5.550 ;
        RECT 13.050 -10.000 13.350 -9.950 ;
        RECT 8.750 -10.400 13.350 -10.000 ;
        RECT 6.350 -10.800 9.150 -10.400 ;
        RECT 13.050 -10.450 13.350 -10.400 ;
        RECT 6.350 -11.145 6.550 -10.800 ;
        RECT 6.315 -11.475 6.565 -11.145 ;
        RECT 13.550 -11.150 13.950 -5.550 ;
        RECT 14.450 -9.550 14.850 -4.500 ;
        RECT 14.150 -10.450 14.450 -9.950 ;
        RECT 17.450 -11.150 17.850 -5.700 ;
        RECT 18.350 -7.700 18.750 -3.500 ;
        RECT 19.250 -7.700 19.650 -5.700 ;
        RECT 21.300 -7.700 21.700 -5.700 ;
        RECT 22.200 -7.700 22.600 -3.500 ;
        RECT 25.800 -4.000 26.200 -3.500 ;
        RECT 25.800 -4.500 26.900 -4.000 ;
        RECT 18.050 -8.600 19.050 -8.100 ;
        RECT 22.000 -8.600 22.850 -8.100 ;
        RECT 13.550 -11.550 17.850 -11.150 ;
        RECT 5.495 -11.645 6.125 -11.565 ;
        RECT 6.725 -11.645 7.705 -11.565 ;
        RECT 5.495 -11.895 7.705 -11.645 ;
        RECT 18.350 -11.950 18.750 -8.600 ;
        RECT 23.100 -10.800 23.500 -5.700 ;
        RECT 25.800 -6.150 26.200 -4.500 ;
        RECT 26.500 -9.600 26.900 -4.500 ;
        RECT 26.900 -10.500 27.200 -10.000 ;
        RECT 27.400 -10.800 27.800 -5.600 ;
        RECT 28.300 -9.600 28.700 -5.600 ;
        RECT 28.000 -10.500 28.300 -10.000 ;
        RECT 29.900 -10.800 30.400 -0.350 ;
        RECT 44.400 -0.325 45.425 -0.075 ;
        RECT 39.685 -2.055 40.015 -1.245 ;
        RECT 39.685 -2.225 40.400 -2.055 ;
        RECT 39.680 -2.400 40.060 -2.395 ;
        RECT 38.100 -2.600 40.060 -2.400 ;
        RECT 38.100 -4.750 38.400 -2.600 ;
        RECT 39.680 -2.635 40.060 -2.600 ;
        RECT 40.230 -2.465 40.400 -2.225 ;
        RECT 40.605 -2.095 40.775 -1.245 ;
        RECT 41.445 -2.095 41.615 -1.245 ;
        RECT 44.400 -1.600 44.650 -0.325 ;
        RECT 40.605 -2.265 41.615 -2.095 ;
        RECT 41.120 -2.400 41.615 -2.265 ;
        RECT 42.350 -1.850 44.650 -1.600 ;
        RECT 45.165 -1.745 45.335 -1.245 ;
        RECT 42.350 -2.400 42.625 -1.850 ;
        RECT 45.165 -1.915 45.830 -1.745 ;
        RECT 40.230 -2.635 40.730 -2.465 ;
        RECT 40.230 -2.805 40.400 -2.635 ;
        RECT 41.120 -2.650 42.625 -2.400 ;
        RECT 41.120 -2.805 41.615 -2.650 ;
        RECT 45.080 -2.735 45.430 -2.085 ;
        RECT 39.765 -2.975 40.400 -2.805 ;
        RECT 40.605 -2.975 41.615 -2.805 ;
        RECT 45.600 -2.905 45.830 -1.915 ;
        RECT 39.765 -3.455 39.935 -2.975 ;
        RECT 40.605 -3.455 40.775 -2.975 ;
        RECT 41.445 -3.455 41.615 -2.975 ;
        RECT 45.165 -3.075 45.830 -2.905 ;
        RECT 45.165 -3.365 45.335 -3.075 ;
        RECT 46.005 -3.365 46.190 -1.245 ;
        RECT 46.865 -1.670 47.115 -1.245 ;
        RECT 47.325 -1.520 48.430 -1.350 ;
        RECT 46.810 -1.800 47.115 -1.670 ;
        RECT 46.360 -2.995 46.640 -2.045 ;
        RECT 46.810 -2.905 46.980 -1.800 ;
        RECT 47.150 -2.585 47.390 -1.990 ;
        RECT 47.560 -2.055 48.090 -1.690 ;
        RECT 47.560 -2.755 47.730 -2.055 ;
        RECT 48.260 -2.135 48.430 -1.520 ;
        RECT 48.940 -1.575 49.190 -1.245 ;
        RECT 49.415 -1.545 50.300 -1.375 ;
        RECT 48.260 -2.225 48.770 -2.135 ;
        RECT 46.810 -3.035 47.035 -2.905 ;
        RECT 47.205 -2.975 47.730 -2.755 ;
        RECT 47.900 -2.395 48.770 -2.225 ;
        RECT 46.865 -3.175 47.035 -3.035 ;
        RECT 47.900 -3.175 48.070 -2.395 ;
        RECT 48.600 -2.465 48.770 -2.395 ;
        RECT 48.280 -2.645 48.480 -2.615 ;
        RECT 48.940 -2.645 49.110 -1.575 ;
        RECT 49.280 -2.465 49.470 -1.745 ;
        RECT 48.280 -2.945 49.110 -2.645 ;
        RECT 49.640 -2.675 49.960 -1.715 ;
        RECT 46.865 -3.345 47.200 -3.175 ;
        RECT 47.395 -3.345 48.070 -3.175 ;
        RECT 48.940 -3.175 49.110 -2.945 ;
        RECT 49.495 -3.005 49.960 -2.675 ;
        RECT 50.130 -2.385 50.300 -1.545 ;
        RECT 51.030 -1.805 51.370 -1.245 ;
        RECT 50.470 -2.180 51.370 -1.805 ;
        RECT 51.180 -2.385 51.370 -2.180 ;
        RECT 51.880 -2.135 52.210 -1.290 ;
        RECT 52.895 -1.995 53.225 -1.265 ;
        RECT 51.880 -2.215 52.290 -2.135 ;
        RECT 52.055 -2.265 52.290 -2.215 ;
        RECT 50.130 -2.715 51.010 -2.385 ;
        RECT 51.180 -2.715 51.930 -2.385 ;
        RECT 50.130 -3.175 50.300 -2.715 ;
        RECT 51.180 -2.885 51.380 -2.715 ;
        RECT 52.100 -2.845 52.290 -2.265 ;
        RECT 52.045 -2.885 52.290 -2.845 ;
        RECT 48.940 -3.345 49.345 -3.175 ;
        RECT 49.515 -3.345 50.300 -3.175 ;
        RECT 51.050 -3.410 51.380 -2.885 ;
        RECT 51.890 -2.970 52.290 -2.885 ;
        RECT 52.955 -2.385 53.225 -1.995 ;
        RECT 53.800 -2.215 54.135 -1.245 ;
        RECT 52.955 -2.715 53.750 -2.385 ;
        RECT 53.920 -2.400 54.135 -2.215 ;
        RECT 53.920 -2.600 56.100 -2.400 ;
        RECT 51.890 -3.405 52.220 -2.970 ;
        RECT 52.955 -3.095 53.155 -2.715 ;
        RECT 53.920 -2.825 54.135 -2.600 ;
        RECT 54.750 -2.750 56.100 -2.600 ;
        RECT 52.895 -3.365 53.155 -3.095 ;
        RECT 53.880 -3.445 54.135 -2.825 ;
        RECT 54.900 -3.350 55.400 -2.950 ;
        RECT 55.700 -4.750 56.100 -2.750 ;
        RECT 38.100 -5.150 56.100 -4.750 ;
        RECT 42.355 -9.545 42.685 -8.745 ;
        RECT 43.195 -9.525 43.525 -8.745 ;
        RECT 46.565 -9.245 46.735 -8.745 ;
        RECT 46.565 -9.415 47.230 -9.245 ;
        RECT 43.195 -9.545 43.960 -9.525 ;
        RECT 42.355 -9.600 43.960 -9.545 ;
        RECT 46.480 -9.600 46.830 -9.585 ;
        RECT 42.355 -9.715 46.830 -9.600 ;
        RECT 41.895 -10.135 43.525 -9.885 ;
        RECT 43.695 -10.000 46.830 -9.715 ;
        RECT 43.695 -10.305 43.960 -10.000 ;
        RECT 46.480 -10.235 46.830 -10.000 ;
        RECT 23.100 -11.300 30.400 -10.800 ;
        RECT 42.355 -10.485 43.960 -10.305 ;
        RECT 47.000 -10.405 47.230 -9.415 ;
        RECT 42.355 -10.955 42.685 -10.485 ;
        RECT 43.195 -10.955 43.525 -10.485 ;
        RECT 45.000 -10.900 45.550 -10.450 ;
        RECT 46.565 -10.575 47.230 -10.405 ;
        RECT 46.565 -10.865 46.735 -10.575 ;
        RECT 47.405 -10.865 47.590 -8.745 ;
        RECT 48.265 -9.170 48.515 -8.745 ;
        RECT 48.725 -9.020 49.830 -8.850 ;
        RECT 48.210 -9.300 48.515 -9.170 ;
        RECT 47.760 -10.495 48.040 -9.545 ;
        RECT 48.210 -10.405 48.380 -9.300 ;
        RECT 48.550 -10.085 48.790 -9.490 ;
        RECT 48.960 -9.555 49.490 -9.190 ;
        RECT 48.960 -10.255 49.130 -9.555 ;
        RECT 49.660 -9.635 49.830 -9.020 ;
        RECT 50.340 -9.075 50.590 -8.745 ;
        RECT 50.815 -9.045 51.700 -8.875 ;
        RECT 49.660 -9.725 50.170 -9.635 ;
        RECT 48.210 -10.535 48.435 -10.405 ;
        RECT 48.605 -10.475 49.130 -10.255 ;
        RECT 49.300 -9.895 50.170 -9.725 ;
        RECT 48.265 -10.675 48.435 -10.535 ;
        RECT 49.300 -10.675 49.470 -9.895 ;
        RECT 50.000 -9.965 50.170 -9.895 ;
        RECT 49.680 -10.145 49.880 -10.115 ;
        RECT 50.340 -10.145 50.510 -9.075 ;
        RECT 50.680 -9.965 50.870 -9.245 ;
        RECT 49.680 -10.445 50.510 -10.145 ;
        RECT 51.040 -10.175 51.360 -9.215 ;
        RECT 48.265 -10.845 48.600 -10.675 ;
        RECT 48.795 -10.845 49.470 -10.675 ;
        RECT 50.340 -10.675 50.510 -10.445 ;
        RECT 50.895 -10.505 51.360 -10.175 ;
        RECT 51.530 -9.885 51.700 -9.045 ;
        RECT 52.425 -9.305 52.765 -8.745 ;
        RECT 51.870 -9.680 52.765 -9.305 ;
        RECT 52.575 -9.885 52.765 -9.680 ;
        RECT 53.275 -9.635 53.605 -8.790 ;
        RECT 53.275 -9.715 53.665 -9.635 ;
        RECT 53.450 -9.765 53.665 -9.715 ;
        RECT 51.530 -10.215 52.405 -9.885 ;
        RECT 52.575 -10.215 53.325 -9.885 ;
        RECT 51.530 -10.675 51.700 -10.215 ;
        RECT 52.575 -10.385 52.775 -10.215 ;
        RECT 53.495 -10.345 53.665 -9.765 ;
        RECT 53.440 -10.385 53.665 -10.345 ;
        RECT 50.340 -10.845 50.745 -10.675 ;
        RECT 50.915 -10.845 51.700 -10.675 ;
        RECT 45.175 -11.775 45.425 -10.900 ;
        RECT 52.445 -10.910 52.775 -10.385 ;
        RECT 53.285 -10.470 53.665 -10.385 ;
        RECT 53.285 -10.905 53.615 -10.470 ;
        RECT 8.750 -12.450 28.700 -11.950 ;
        RECT 44.400 -12.025 45.425 -11.775 ;
        RECT 8.750 -13.050 9.250 -12.450 ;
        RECT 6.600 -13.550 9.250 -13.050 ;
        RECT 39.685 -13.755 40.015 -12.945 ;
        RECT 39.685 -13.925 40.400 -13.755 ;
        RECT 39.680 -14.100 40.060 -14.095 ;
        RECT 38.100 -14.300 40.060 -14.100 ;
        RECT 14.830 -15.270 16.990 -14.920 ;
        RECT 38.100 -16.450 38.400 -14.300 ;
        RECT 39.680 -14.335 40.060 -14.300 ;
        RECT 40.230 -14.165 40.400 -13.925 ;
        RECT 40.605 -13.795 40.775 -12.945 ;
        RECT 41.445 -13.795 41.615 -12.945 ;
        RECT 44.400 -13.300 44.650 -12.025 ;
        RECT 40.605 -13.965 41.615 -13.795 ;
        RECT 41.120 -14.100 41.615 -13.965 ;
        RECT 42.350 -13.550 44.650 -13.300 ;
        RECT 45.165 -13.445 45.335 -12.945 ;
        RECT 42.350 -14.100 42.625 -13.550 ;
        RECT 45.165 -13.615 45.830 -13.445 ;
        RECT 40.230 -14.335 40.730 -14.165 ;
        RECT 40.230 -14.505 40.400 -14.335 ;
        RECT 41.120 -14.350 42.625 -14.100 ;
        RECT 41.120 -14.505 41.615 -14.350 ;
        RECT 45.080 -14.435 45.430 -13.785 ;
        RECT 39.765 -14.675 40.400 -14.505 ;
        RECT 40.605 -14.675 41.615 -14.505 ;
        RECT 45.600 -14.605 45.830 -13.615 ;
        RECT 39.765 -15.155 39.935 -14.675 ;
        RECT 40.605 -15.155 40.775 -14.675 ;
        RECT 41.445 -15.155 41.615 -14.675 ;
        RECT 45.165 -14.775 45.830 -14.605 ;
        RECT 45.165 -15.065 45.335 -14.775 ;
        RECT 46.005 -15.065 46.190 -12.945 ;
        RECT 46.865 -13.370 47.115 -12.945 ;
        RECT 47.325 -13.220 48.430 -13.050 ;
        RECT 46.810 -13.500 47.115 -13.370 ;
        RECT 46.360 -14.695 46.640 -13.745 ;
        RECT 46.810 -14.605 46.980 -13.500 ;
        RECT 47.150 -14.285 47.390 -13.690 ;
        RECT 47.560 -13.755 48.090 -13.390 ;
        RECT 47.560 -14.455 47.730 -13.755 ;
        RECT 48.260 -13.835 48.430 -13.220 ;
        RECT 48.940 -13.275 49.190 -12.945 ;
        RECT 49.415 -13.245 50.300 -13.075 ;
        RECT 48.260 -13.925 48.770 -13.835 ;
        RECT 46.810 -14.735 47.035 -14.605 ;
        RECT 47.205 -14.675 47.730 -14.455 ;
        RECT 47.900 -14.095 48.770 -13.925 ;
        RECT 46.865 -14.875 47.035 -14.735 ;
        RECT 47.900 -14.875 48.070 -14.095 ;
        RECT 48.600 -14.165 48.770 -14.095 ;
        RECT 48.280 -14.345 48.480 -14.315 ;
        RECT 48.940 -14.345 49.110 -13.275 ;
        RECT 49.280 -14.165 49.470 -13.445 ;
        RECT 48.280 -14.645 49.110 -14.345 ;
        RECT 49.640 -14.375 49.960 -13.415 ;
        RECT 46.865 -15.045 47.200 -14.875 ;
        RECT 47.395 -15.045 48.070 -14.875 ;
        RECT 48.940 -14.875 49.110 -14.645 ;
        RECT 49.495 -14.705 49.960 -14.375 ;
        RECT 50.130 -14.085 50.300 -13.245 ;
        RECT 51.030 -13.505 51.370 -12.945 ;
        RECT 50.470 -13.880 51.370 -13.505 ;
        RECT 52.895 -13.695 53.225 -12.965 ;
        RECT 51.180 -14.085 51.370 -13.880 ;
        RECT 52.955 -14.085 53.225 -13.695 ;
        RECT 53.800 -13.915 54.135 -12.945 ;
        RECT 50.130 -14.415 51.010 -14.085 ;
        RECT 51.180 -14.415 51.930 -14.085 ;
        RECT 52.955 -14.415 53.750 -14.085 ;
        RECT 53.920 -14.100 54.135 -13.915 ;
        RECT 53.920 -14.300 56.100 -14.100 ;
        RECT 50.130 -14.875 50.300 -14.415 ;
        RECT 51.180 -14.585 51.380 -14.415 ;
        RECT 48.940 -15.045 49.345 -14.875 ;
        RECT 49.515 -15.045 50.300 -14.875 ;
        RECT 51.050 -15.110 51.380 -14.585 ;
        RECT 52.955 -14.795 53.155 -14.415 ;
        RECT 53.920 -14.525 54.135 -14.300 ;
        RECT 54.750 -14.450 56.100 -14.300 ;
        RECT 52.895 -15.065 53.155 -14.795 ;
        RECT 53.880 -15.145 54.135 -14.525 ;
        RECT 54.900 -15.050 55.400 -14.650 ;
        RECT 55.700 -16.450 56.100 -14.450 ;
        RECT 38.100 -16.850 56.100 -16.450 ;
      LAYER met1 ;
        RECT 8.600 30.400 55.600 30.800 ;
        RECT 8.600 27.850 9.000 30.400 ;
        RECT 12.900 27.750 13.300 30.400 ;
        RECT 15.800 27.750 16.200 30.400 ;
        RECT 18.700 27.850 19.100 30.400 ;
        RECT 23.000 27.850 23.400 30.400 ;
        RECT 27.300 27.750 27.700 30.400 ;
        RECT 30.200 27.750 30.600 30.400 ;
        RECT 33.100 27.850 33.500 30.400 ;
        RECT 37.400 27.850 37.800 30.400 ;
        RECT 41.700 27.750 42.100 30.400 ;
        RECT 44.600 27.750 45.000 30.400 ;
        RECT 47.500 27.850 47.900 30.400 ;
        RECT 10.700 27.300 11.100 27.500 ;
        RECT 17.900 27.300 18.300 27.500 ;
        RECT 10.700 27.100 18.300 27.300 ;
        RECT 25.100 27.300 25.500 27.500 ;
        RECT 32.300 27.300 32.700 27.500 ;
        RECT 25.100 27.100 32.700 27.300 ;
        RECT 39.500 27.300 39.900 27.500 ;
        RECT 46.700 27.300 47.100 27.500 ;
        RECT 39.500 27.100 47.100 27.300 ;
        RECT 5.900 26.700 10.350 27.100 ;
        RECT 10.700 26.900 24.750 27.100 ;
        RECT 10.700 26.700 11.100 26.900 ;
        RECT 5.900 11.500 6.400 26.700 ;
        RECT 9.950 24.950 10.350 26.700 ;
        RECT 9.950 24.500 11.800 24.950 ;
        RECT 14.250 24.550 14.650 26.900 ;
        RECT 17.900 26.700 24.750 26.900 ;
        RECT 25.100 26.900 39.150 27.100 ;
        RECT 25.100 26.700 25.500 26.900 ;
        RECT 17.900 26.300 18.300 26.700 ;
        RECT 15.000 25.500 21.200 25.900 ;
        RECT 17.150 24.550 17.550 25.500 ;
        RECT 24.350 24.950 24.750 26.700 ;
        RECT 20.050 24.500 21.900 24.950 ;
        RECT 24.350 24.500 26.200 24.950 ;
        RECT 28.650 24.550 29.050 26.900 ;
        RECT 32.300 26.700 39.150 26.900 ;
        RECT 39.500 26.900 54.100 27.100 ;
        RECT 39.500 26.700 39.900 26.900 ;
        RECT 32.300 26.300 32.700 26.700 ;
        RECT 29.400 25.500 35.600 25.900 ;
        RECT 31.550 24.550 31.950 25.500 ;
        RECT 38.750 24.950 39.150 26.700 ;
        RECT 34.450 24.500 36.300 24.950 ;
        RECT 38.750 24.500 40.600 24.950 ;
        RECT 43.050 24.550 43.450 26.900 ;
        RECT 46.700 26.700 54.100 26.900 ;
        RECT 46.700 26.300 47.100 26.700 ;
        RECT 43.800 25.500 50.000 25.900 ;
        RECT 45.950 24.550 46.350 25.500 ;
        RECT 48.850 24.500 50.700 24.950 ;
        RECT 20.050 23.400 20.500 24.500 ;
        RECT 7.400 23.000 20.500 23.400 ;
        RECT 20.800 23.400 21.200 23.800 ;
        RECT 34.450 23.400 34.900 24.500 ;
        RECT 20.800 23.000 34.900 23.400 ;
        RECT 35.200 23.400 35.600 23.800 ;
        RECT 48.850 23.400 49.300 24.500 ;
        RECT 35.200 23.000 49.300 23.400 ;
        RECT 49.600 23.400 50.000 23.800 ;
        RECT 49.600 23.000 52.600 23.400 ;
        RECT 7.400 15.200 7.900 23.000 ;
        RECT 20.800 22.600 21.200 23.000 ;
        RECT 35.200 22.600 35.600 23.000 ;
        RECT 49.600 22.600 50.000 23.000 ;
        RECT 24.450 15.200 24.850 15.600 ;
        RECT 38.850 15.200 39.250 15.600 ;
        RECT 52.100 15.200 52.600 23.000 ;
        RECT 7.400 14.800 24.850 15.200 ;
        RECT 24.450 14.400 24.850 14.800 ;
        RECT 25.150 14.800 39.250 15.200 ;
        RECT 25.150 13.700 25.600 14.800 ;
        RECT 38.850 14.400 39.250 14.800 ;
        RECT 39.550 14.800 52.600 15.200 ;
        RECT 39.550 13.700 40.000 14.800 ;
        RECT 23.750 13.250 25.600 13.700 ;
        RECT 28.100 12.700 28.500 13.650 ;
        RECT 24.450 12.300 30.650 12.700 ;
        RECT 27.350 11.500 27.750 11.900 ;
        RECT 5.900 11.300 27.750 11.500 ;
        RECT 31.000 11.300 31.400 13.650 ;
        RECT 33.850 13.250 35.700 13.700 ;
        RECT 38.150 13.250 40.000 13.700 ;
        RECT 35.300 11.500 35.700 13.250 ;
        RECT 42.500 12.700 42.900 13.650 ;
        RECT 38.850 12.300 45.050 12.700 ;
        RECT 41.750 11.500 42.150 11.900 ;
        RECT 34.550 11.300 34.950 11.500 ;
        RECT 5.900 11.100 34.950 11.300 ;
        RECT 35.300 11.300 42.150 11.500 ;
        RECT 45.400 11.300 45.800 13.650 ;
        RECT 48.250 13.250 50.100 13.700 ;
        RECT 49.700 11.500 50.100 13.250 ;
        RECT 53.600 11.500 54.100 26.700 ;
        RECT 48.950 11.300 49.350 11.500 ;
        RECT 35.300 11.100 49.350 11.300 ;
        RECT 49.700 11.100 54.100 11.500 ;
        RECT 21.100 6.200 21.500 11.100 ;
        RECT 27.350 10.900 34.950 11.100 ;
        RECT 27.350 10.700 27.750 10.900 ;
        RECT 34.550 10.700 34.950 10.900 ;
        RECT 41.750 10.900 49.350 11.100 ;
        RECT 41.750 10.700 42.150 10.900 ;
        RECT 48.950 10.700 49.350 10.900 ;
        RECT 26.550 7.800 26.950 10.350 ;
        RECT 29.450 7.800 29.850 10.450 ;
        RECT 32.350 7.800 32.750 10.450 ;
        RECT 36.650 7.800 37.050 10.350 ;
        RECT 40.950 7.800 41.350 10.350 ;
        RECT 43.850 7.800 44.250 10.450 ;
        RECT 46.750 7.800 47.150 10.450 ;
        RECT 51.050 7.800 51.450 10.350 ;
        RECT 55.100 7.800 55.600 30.400 ;
        RECT 26.550 7.400 55.600 7.800 ;
        RECT 21.100 5.800 32.450 6.200 ;
        RECT 32.050 4.550 32.450 5.800 ;
        RECT 32.050 4.540 34.150 4.550 ;
        RECT 32.050 4.180 34.480 4.540 ;
        RECT 35.100 4.500 35.350 5.500 ;
        RECT 36.750 4.500 41.350 4.650 ;
        RECT 35.100 4.300 41.350 4.500 ;
        RECT 35.185 4.290 41.350 4.300 ;
        RECT 32.050 4.150 34.150 4.180 ;
        RECT 36.750 4.150 41.350 4.290 ;
        RECT 40.850 1.900 41.350 4.150 ;
        RECT 46.960 2.430 47.250 2.475 ;
        RECT 49.060 2.430 49.350 2.475 ;
        RECT 50.630 2.430 50.920 2.475 ;
        RECT 46.960 2.290 50.920 2.430 ;
        RECT 46.960 2.245 47.250 2.290 ;
        RECT 49.060 2.245 49.350 2.290 ;
        RECT 50.630 2.245 50.920 2.290 ;
        RECT 47.355 2.090 47.645 2.135 ;
        RECT 48.545 2.090 48.835 2.135 ;
        RECT 51.065 2.090 51.355 2.135 ;
        RECT 47.355 1.950 51.355 2.090 ;
        RECT 47.355 1.905 47.645 1.950 ;
        RECT 48.545 1.905 48.835 1.950 ;
        RECT 51.065 1.905 51.355 1.950 ;
        RECT 39.100 1.600 42.300 1.900 ;
        RECT 20.850 1.050 21.250 1.550 ;
        RECT 21.550 1.400 21.950 1.500 ;
        RECT 23.350 1.400 23.750 1.500 ;
        RECT 21.550 0.850 23.750 1.400 ;
        RECT 21.550 0.700 21.950 0.850 ;
        RECT 23.350 0.700 23.750 0.850 ;
        RECT 13.200 -2.200 13.600 0.700 ;
        RECT 16.950 -0.200 19.150 0.300 ;
        RECT 16.950 -0.300 17.350 -0.200 ;
        RECT 18.750 -0.300 19.150 -0.200 ;
        RECT 22.450 -0.300 24.650 0.300 ;
        RECT 26.350 -2.200 26.750 1.500 ;
        RECT 27.050 -2.200 27.450 0.650 ;
        RECT 39.100 -0.100 39.400 1.600 ;
        RECT 41.900 1.500 42.300 1.600 ;
        RECT 47.650 1.350 48.150 1.700 ;
        RECT 45.000 1.000 48.150 1.350 ;
        RECT 45.000 0.800 45.550 1.000 ;
        RECT 53.300 0.900 58.250 1.400 ;
        RECT 39.100 -0.400 43.050 -0.100 ;
        RECT 13.200 -2.600 27.450 -2.200 ;
        RECT 42.750 -2.450 43.050 -0.400 ;
        RECT 55.400 -1.400 55.900 -0.250 ;
        RECT 51.850 -1.650 55.900 -1.400 ;
        RECT 45.560 -1.770 45.850 -1.725 ;
        RECT 47.660 -1.770 47.950 -1.725 ;
        RECT 49.230 -1.770 49.520 -1.725 ;
        RECT 45.560 -1.910 49.520 -1.770 ;
        RECT 45.560 -1.955 45.850 -1.910 ;
        RECT 47.660 -1.955 47.950 -1.910 ;
        RECT 49.230 -1.955 49.520 -1.910 ;
        RECT 45.050 -2.450 45.450 -2.100 ;
        RECT 45.955 -2.110 46.245 -2.065 ;
        RECT 47.145 -2.110 47.435 -2.065 ;
        RECT 49.665 -2.110 49.955 -2.065 ;
        RECT 45.955 -2.250 49.955 -2.110 ;
        RECT 45.955 -2.295 46.245 -2.250 ;
        RECT 47.145 -2.295 47.435 -2.250 ;
        RECT 49.665 -2.295 49.955 -2.250 ;
        RECT 42.750 -2.750 45.450 -2.450 ;
        RECT 46.350 -3.000 46.750 -2.400 ;
        RECT 44.000 -3.250 46.750 -3.000 ;
        RECT 51.850 -2.450 52.300 -1.650 ;
        RECT 51.850 -3.200 52.350 -2.450 ;
        RECT 15.450 -4.950 20.850 -4.450 ;
        RECT 11.950 -6.000 12.350 -5.500 ;
        RECT 12.650 -5.700 13.050 -5.550 ;
        RECT 14.450 -5.700 14.850 -5.550 ;
        RECT 12.650 -6.200 14.850 -5.700 ;
        RECT 12.650 -6.350 13.050 -6.200 ;
        RECT 14.450 -6.350 14.850 -6.200 ;
        RECT 12.650 -8.900 13.050 -8.750 ;
        RECT 14.450 -8.900 14.850 -8.750 ;
        RECT 12.650 -9.400 14.850 -8.900 ;
        RECT 12.650 -9.550 13.050 -9.400 ;
        RECT 14.450 -9.550 14.850 -9.400 ;
        RECT 15.450 -9.950 15.950 -4.950 ;
        RECT 17.450 -5.900 17.850 -5.700 ;
        RECT 19.250 -5.900 19.650 -5.700 ;
        RECT 17.450 -6.400 19.650 -5.900 ;
        RECT 17.450 -6.550 17.850 -6.400 ;
        RECT 19.250 -6.550 19.650 -6.400 ;
        RECT 20.350 -8.100 20.850 -4.950 ;
        RECT 44.000 -5.500 44.500 -3.250 ;
        RECT 54.900 -3.350 55.400 -2.950 ;
        RECT 57.750 -5.500 58.250 0.900 ;
        RECT 21.300 -6.200 21.700 -5.700 ;
        RECT 23.100 -6.200 23.500 -5.700 ;
        RECT 25.800 -6.150 26.200 -5.650 ;
        RECT 26.500 -5.750 26.900 -5.600 ;
        RECT 28.300 -5.750 28.700 -5.600 ;
        RECT 21.300 -6.700 23.500 -6.200 ;
        RECT 26.500 -6.250 28.700 -5.750 ;
        RECT 44.000 -6.000 58.250 -5.500 ;
        RECT 26.500 -6.400 26.900 -6.250 ;
        RECT 28.300 -6.400 28.700 -6.250 ;
        RECT 21.300 -6.850 21.700 -6.700 ;
        RECT 23.100 -6.850 23.500 -6.700 ;
        RECT 59.200 -7.150 59.700 -0.250 ;
        RECT 40.700 -7.650 59.700 -7.150 ;
        RECT 17.850 -8.600 19.250 -8.100 ;
        RECT 20.350 -8.600 23.100 -8.100 ;
        RECT 26.500 -8.950 26.900 -8.800 ;
        RECT 28.300 -8.950 28.700 -8.800 ;
        RECT 26.500 -9.450 28.700 -8.950 ;
        RECT 26.500 -9.600 26.900 -9.450 ;
        RECT 28.300 -9.600 28.700 -9.450 ;
        RECT 40.700 -9.800 41.200 -7.650 ;
        RECT 46.960 -9.270 47.250 -9.225 ;
        RECT 49.060 -9.270 49.350 -9.225 ;
        RECT 50.630 -9.270 50.920 -9.225 ;
        RECT 46.960 -9.410 50.920 -9.270 ;
        RECT 46.960 -9.455 47.250 -9.410 ;
        RECT 49.060 -9.455 49.350 -9.410 ;
        RECT 50.630 -9.455 50.920 -9.410 ;
        RECT 47.355 -9.610 47.645 -9.565 ;
        RECT 48.545 -9.610 48.835 -9.565 ;
        RECT 51.065 -9.610 51.355 -9.565 ;
        RECT 47.355 -9.750 51.355 -9.610 ;
        RECT 47.355 -9.795 47.645 -9.750 ;
        RECT 48.545 -9.795 48.835 -9.750 ;
        RECT 51.065 -9.795 51.355 -9.750 ;
        RECT 13.050 -10.450 15.950 -9.950 ;
        RECT 26.900 -10.500 28.700 -10.000 ;
        RECT 6.600 -11.900 7.450 -11.550 ;
        RECT 13.350 -11.700 14.150 -11.000 ;
        RECT 6.600 -13.550 7.100 -11.900 ;
        RECT 13.550 -14.900 13.950 -11.700 ;
        RECT 28.300 -12.450 28.700 -10.500 ;
        RECT 39.100 -10.100 42.300 -9.800 ;
        RECT 39.100 -11.800 39.400 -10.100 ;
        RECT 41.900 -10.200 42.300 -10.100 ;
        RECT 47.650 -10.350 48.150 -10.000 ;
        RECT 45.000 -10.700 48.150 -10.350 ;
        RECT 45.000 -10.900 45.550 -10.700 ;
        RECT 53.300 -10.800 58.250 -10.300 ;
        RECT 39.100 -12.100 43.050 -11.800 ;
        RECT 42.750 -14.150 43.050 -12.100 ;
        RECT 45.560 -13.470 45.850 -13.425 ;
        RECT 47.660 -13.470 47.950 -13.425 ;
        RECT 49.230 -13.470 49.520 -13.425 ;
        RECT 45.560 -13.610 49.520 -13.470 ;
        RECT 45.560 -13.655 45.850 -13.610 ;
        RECT 47.660 -13.655 47.950 -13.610 ;
        RECT 49.230 -13.655 49.520 -13.610 ;
        RECT 45.050 -14.150 45.450 -13.800 ;
        RECT 45.955 -13.810 46.245 -13.765 ;
        RECT 47.145 -13.810 47.435 -13.765 ;
        RECT 49.665 -13.810 49.955 -13.765 ;
        RECT 45.955 -13.950 49.955 -13.810 ;
        RECT 45.955 -13.995 46.245 -13.950 ;
        RECT 47.145 -13.995 47.435 -13.950 ;
        RECT 49.665 -13.995 49.955 -13.950 ;
        RECT 42.750 -14.450 45.450 -14.150 ;
        RECT 46.350 -14.700 46.750 -14.100 ;
        RECT 13.550 -14.970 15.000 -14.900 ;
        RECT 44.000 -14.950 46.750 -14.700 ;
        RECT 13.550 -15.220 16.965 -14.970 ;
        RECT 13.550 -15.300 15.000 -15.220 ;
        RECT 44.000 -17.200 44.500 -14.950 ;
        RECT 54.900 -15.050 55.400 -14.650 ;
        RECT 57.750 -17.200 58.250 -10.800 ;
        RECT 44.000 -17.700 58.250 -17.200 ;
      LAYER met2 ;
        RECT 55.400 -0.750 59.700 -0.250 ;
  END
END dco
MACRO qz
  CLASS BLOCK ;
  FOREIGN qz ;
  ORIGIN -0.950 3.550 ;
  SIZE 28.500 BY 7.200 ;
  PIN CLK
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.745 4.415 2.305 ;
        RECT 7.530 -2.335 7.880 -1.685 ;
      LAYER met1 ;
        RECT 3.730 2.200 4.430 2.320 ;
        RECT 2.200 1.850 4.430 2.200 ;
        RECT 2.200 0.200 2.550 1.850 ;
        RECT 3.730 1.750 4.430 1.850 ;
        RECT 2.200 -0.150 7.050 0.200 ;
        RECT 6.700 -1.650 7.050 -0.150 ;
        RECT 6.700 -1.690 7.850 -1.650 ;
        RECT 6.700 -2.000 7.860 -1.690 ;
        RECT 7.510 -2.340 7.860 -2.000 ;
    END
  END CLK
  PIN Dout
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 14.325 -1.735 14.655 -0.890 ;
        RECT 14.325 -1.815 14.715 -1.735 ;
        RECT 14.500 -1.865 14.715 -1.815 ;
        RECT 14.545 -2.000 14.715 -1.865 ;
        RECT 16.785 -2.000 17.120 -1.985 ;
        RECT 14.545 -2.250 17.120 -2.000 ;
        RECT 14.545 -2.445 14.715 -2.250 ;
        RECT 16.785 -2.255 17.120 -2.250 ;
        RECT 14.490 -2.485 14.715 -2.445 ;
        RECT 14.335 -2.570 14.715 -2.485 ;
        RECT 14.335 -3.005 14.665 -2.570 ;
    END
  END Dout
  PIN FBack
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 19.865 -1.825 20.195 -0.845 ;
        RECT 19.945 -2.425 20.195 -1.825 ;
        RECT 19.865 -3.055 20.195 -2.425 ;
      LAYER met1 ;
        RECT 19.850 -1.250 20.250 -1.100 ;
        RECT 19.850 -1.600 21.850 -1.250 ;
    END
  END FBack
  PIN D
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.725 -2.325 4.080 -1.955 ;
      LAYER met1 ;
        RECT 3.700 -1.950 4.100 -1.900 ;
        RECT 2.200 -2.300 4.100 -1.950 ;
        RECT 3.700 -2.350 4.100 -2.300 ;
    END
  END D
  PIN GND
    ANTENNADIFFAREA 3.821850 ;
    PORT
      LAYER pwell ;
        RECT 3.450 0.750 28.350 1.750 ;
        RECT 3.785 0.605 3.955 0.750 ;
        RECT 7.885 0.605 8.055 0.750 ;
        RECT 11.985 0.605 12.155 0.750 ;
        RECT 16.385 0.605 16.555 0.750 ;
        RECT 20.485 0.605 20.655 0.750 ;
        RECT 24.585 0.605 24.755 0.750 ;
        RECT 3.450 -3.250 20.950 -2.250 ;
        RECT 3.785 -3.395 3.955 -3.250 ;
        RECT 7.585 -3.395 7.755 -3.250 ;
        RECT 16.830 -3.395 17.000 -3.250 ;
        RECT 19.485 -3.395 19.655 -3.250 ;
      LAYER li1 ;
        RECT 4.295 0.775 4.565 1.235 ;
        RECT 6.355 0.775 6.680 1.235 ;
        RECT 8.395 0.775 8.665 1.235 ;
        RECT 10.455 0.775 10.780 1.235 ;
        RECT 12.495 0.775 12.765 1.235 ;
        RECT 14.555 0.775 14.880 1.235 ;
        RECT 15.700 0.940 16.010 1.440 ;
        RECT 16.895 0.775 17.165 1.235 ;
        RECT 18.955 0.775 19.280 1.235 ;
        RECT 20.995 0.775 21.265 1.235 ;
        RECT 23.055 0.775 23.380 1.235 ;
        RECT 25.095 0.775 25.365 1.235 ;
        RECT 27.155 0.775 27.480 1.235 ;
        RECT 3.640 0.605 7.320 0.775 ;
        RECT 7.740 0.605 11.420 0.775 ;
        RECT 11.840 0.605 15.520 0.775 ;
        RECT 16.240 0.605 19.920 0.775 ;
        RECT 20.340 0.605 24.020 0.775 ;
        RECT 24.440 0.605 28.120 0.775 ;
        RECT 4.200 -3.225 4.530 -2.845 ;
        RECT 5.130 -3.225 5.390 -2.385 ;
        RECT 5.650 -2.950 6.050 -2.450 ;
        RECT 7.955 -3.225 8.285 -2.845 ;
        RECT 8.895 -3.225 9.145 -2.765 ;
        RECT 10.840 -3.225 11.210 -2.725 ;
        RECT 13.025 -3.225 13.235 -2.695 ;
        RECT 13.995 -3.225 14.165 -2.615 ;
        RECT 16.775 -3.225 17.085 -2.425 ;
        RECT 19.465 -3.225 19.695 -2.405 ;
        RECT 20.365 -3.225 20.575 -2.405 ;
        RECT 3.640 -3.395 5.480 -3.225 ;
        RECT 7.440 -3.395 14.800 -3.225 ;
        RECT 16.690 -3.395 18.070 -3.225 ;
        RECT 19.340 -3.395 20.720 -3.225 ;
      LAYER met1 ;
        RECT 15.700 0.950 16.010 1.440 ;
        RECT 7.300 0.930 7.750 0.950 ;
        RECT 11.400 0.930 11.850 0.950 ;
        RECT 15.500 0.930 16.250 0.950 ;
        RECT 19.900 0.930 20.350 0.950 ;
        RECT 24.000 0.930 24.450 0.950 ;
        RECT 3.640 0.450 28.120 0.930 ;
        RECT 5.650 -3.050 6.050 -2.450 ;
        RECT 23.460 -3.050 23.935 0.450 ;
        RECT 5.450 -3.070 7.450 -3.050 ;
        RECT 14.800 -3.070 16.700 -3.050 ;
        RECT 18.050 -3.070 19.350 -3.050 ;
        RECT 20.650 -3.070 23.935 -3.050 ;
        RECT 3.640 -3.550 23.935 -3.070 ;
    END
  END GND
  PIN VCCD
    ANTENNADIFFAREA 5.393450 ;
    PORT
      LAYER nwell ;
        RECT 3.650 3.600 28.350 3.650 ;
        RECT 3.450 1.950 28.350 3.600 ;
        RECT 4.600 -0.400 20.950 -0.350 ;
        RECT 3.450 -2.050 20.950 -0.400 ;
      LAYER li1 ;
        RECT 3.650 3.495 4.050 3.650 ;
        RECT 3.640 3.325 7.320 3.495 ;
        RECT 7.740 3.325 11.420 3.495 ;
        RECT 11.840 3.325 15.520 3.495 ;
        RECT 16.240 3.325 19.920 3.495 ;
        RECT 20.340 3.325 24.020 3.495 ;
        RECT 24.440 3.325 28.120 3.495 ;
        RECT 4.295 2.865 4.565 3.325 ;
        RECT 6.355 2.865 6.680 3.325 ;
        RECT 8.395 2.865 8.665 3.325 ;
        RECT 10.455 2.865 10.780 3.325 ;
        RECT 12.495 2.865 12.765 3.325 ;
        RECT 14.555 2.865 14.880 3.325 ;
        RECT 15.750 2.500 16.150 3.000 ;
        RECT 16.895 2.865 17.165 3.325 ;
        RECT 18.955 2.865 19.280 3.325 ;
        RECT 20.995 2.865 21.265 3.325 ;
        RECT 23.055 2.865 23.380 3.325 ;
        RECT 25.095 2.865 25.365 3.325 ;
        RECT 27.155 2.865 27.480 3.325 ;
        RECT 5.100 -0.505 7.850 -0.350 ;
        RECT 3.640 -0.550 14.800 -0.505 ;
        RECT 3.640 -0.675 5.480 -0.550 ;
        RECT 4.200 -1.435 4.530 -0.675 ;
        RECT 5.130 -1.825 5.390 -0.675 ;
        RECT 5.900 -1.500 6.300 -0.550 ;
        RECT 7.440 -0.675 14.800 -0.550 ;
        RECT 16.690 -0.675 18.070 -0.505 ;
        RECT 19.340 -0.675 20.720 -0.505 ;
        RECT 7.955 -1.175 8.285 -0.675 ;
        RECT 8.880 -1.135 9.145 -0.675 ;
        RECT 11.050 -1.475 11.220 -0.675 ;
        RECT 12.930 -1.175 13.245 -0.675 ;
        RECT 13.985 -1.685 14.155 -0.675 ;
        RECT 16.775 -1.815 17.055 -0.675 ;
        RECT 17.725 -1.815 17.985 -0.675 ;
        RECT 19.465 -1.815 19.695 -0.675 ;
        RECT 20.365 -1.815 20.575 -0.675 ;
      LAYER met1 ;
        RECT 0.950 3.170 28.120 3.650 ;
        RECT 0.950 3.150 3.750 3.170 ;
        RECT 7.300 3.150 7.800 3.170 ;
        RECT 11.400 3.150 11.900 3.170 ;
        RECT 15.500 3.150 16.250 3.170 ;
        RECT 19.900 3.150 20.350 3.170 ;
        RECT 24.000 3.150 24.450 3.170 ;
        RECT 0.950 -0.350 1.450 3.150 ;
        RECT 15.750 2.500 16.150 3.150 ;
        RECT 0.950 -0.830 5.480 -0.350 ;
        RECT 7.440 -0.830 20.720 -0.350 ;
        RECT 0.950 -0.850 3.750 -0.830 ;
        RECT 14.800 -0.850 16.700 -0.830 ;
        RECT 18.050 -0.850 19.350 -0.830 ;
        RECT 5.900 -1.500 6.300 -1.000 ;
    END
  END VCCD
  OBS
      LAYER li1 ;
        RECT 3.840 2.695 4.125 3.155 ;
        RECT 3.840 2.475 4.795 2.695 ;
        RECT 4.585 1.575 4.795 2.475 ;
        RECT 3.840 1.405 4.795 1.575 ;
        RECT 4.965 2.305 5.365 3.155 ;
        RECT 5.555 2.695 5.835 3.155 ;
        RECT 5.555 2.475 6.680 2.695 ;
        RECT 4.965 1.745 6.060 2.305 ;
        RECT 6.230 2.015 6.680 2.475 ;
        RECT 6.850 2.300 7.235 3.155 ;
        RECT 7.940 2.695 8.225 3.155 ;
        RECT 7.940 2.475 8.895 2.695 ;
        RECT 7.825 2.300 8.515 2.305 ;
        RECT 6.850 2.185 8.515 2.300 ;
        RECT 3.840 0.945 4.125 1.405 ;
        RECT 4.965 0.945 5.365 1.745 ;
        RECT 6.230 1.685 6.785 2.015 ;
        RECT 6.955 1.750 8.515 2.185 ;
        RECT 6.230 1.575 6.680 1.685 ;
        RECT 5.555 1.405 6.680 1.575 ;
        RECT 6.955 1.515 7.235 1.750 ;
        RECT 7.825 1.745 8.515 1.750 ;
        RECT 8.685 1.575 8.895 2.475 ;
        RECT 5.555 0.945 5.835 1.405 ;
        RECT 6.850 0.945 7.235 1.515 ;
        RECT 7.940 1.405 8.895 1.575 ;
        RECT 9.065 2.305 9.465 3.155 ;
        RECT 9.655 2.695 9.935 3.155 ;
        RECT 9.655 2.475 10.780 2.695 ;
        RECT 9.065 1.745 10.160 2.305 ;
        RECT 10.330 2.015 10.780 2.475 ;
        RECT 10.950 2.300 11.335 3.155 ;
        RECT 12.040 2.695 12.325 3.155 ;
        RECT 12.040 2.475 12.995 2.695 ;
        RECT 11.925 2.300 12.615 2.305 ;
        RECT 10.950 2.185 12.615 2.300 ;
        RECT 7.940 0.945 8.225 1.405 ;
        RECT 9.065 0.945 9.465 1.745 ;
        RECT 10.330 1.685 10.885 2.015 ;
        RECT 11.055 1.750 12.615 2.185 ;
        RECT 10.330 1.575 10.780 1.685 ;
        RECT 9.655 1.405 10.780 1.575 ;
        RECT 11.055 1.515 11.335 1.750 ;
        RECT 11.925 1.745 12.615 1.750 ;
        RECT 12.785 1.575 12.995 2.475 ;
        RECT 9.655 0.945 9.935 1.405 ;
        RECT 10.950 0.945 11.335 1.515 ;
        RECT 12.040 1.405 12.995 1.575 ;
        RECT 13.165 2.305 13.565 3.155 ;
        RECT 13.755 2.695 14.035 3.155 ;
        RECT 13.755 2.475 14.880 2.695 ;
        RECT 13.165 1.745 14.260 2.305 ;
        RECT 14.430 2.015 14.880 2.475 ;
        RECT 15.050 2.300 15.435 3.155 ;
        RECT 16.440 2.695 16.725 3.155 ;
        RECT 16.440 2.475 17.395 2.695 ;
        RECT 16.325 2.300 17.015 2.305 ;
        RECT 15.050 2.185 17.015 2.300 ;
        RECT 12.040 0.945 12.325 1.405 ;
        RECT 13.165 0.945 13.565 1.745 ;
        RECT 14.430 1.685 14.985 2.015 ;
        RECT 15.155 1.750 17.015 2.185 ;
        RECT 14.430 1.575 14.880 1.685 ;
        RECT 13.755 1.405 14.880 1.575 ;
        RECT 15.155 1.515 15.435 1.750 ;
        RECT 16.325 1.745 17.015 1.750 ;
        RECT 17.185 1.575 17.395 2.475 ;
        RECT 13.755 0.945 14.035 1.405 ;
        RECT 15.050 0.945 15.435 1.515 ;
        RECT 16.440 1.405 17.395 1.575 ;
        RECT 17.565 2.305 17.965 3.155 ;
        RECT 18.155 2.695 18.435 3.155 ;
        RECT 18.155 2.475 19.280 2.695 ;
        RECT 17.565 1.745 18.660 2.305 ;
        RECT 18.830 2.015 19.280 2.475 ;
        RECT 19.450 2.300 19.835 3.155 ;
        RECT 20.540 2.695 20.825 3.155 ;
        RECT 20.540 2.475 21.495 2.695 ;
        RECT 20.425 2.300 21.115 2.305 ;
        RECT 19.450 2.185 21.115 2.300 ;
        RECT 16.440 0.945 16.725 1.405 ;
        RECT 17.565 0.945 17.965 1.745 ;
        RECT 18.830 1.685 19.385 2.015 ;
        RECT 19.555 1.750 21.115 2.185 ;
        RECT 18.830 1.575 19.280 1.685 ;
        RECT 18.155 1.405 19.280 1.575 ;
        RECT 19.555 1.515 19.835 1.750 ;
        RECT 20.425 1.745 21.115 1.750 ;
        RECT 21.285 1.575 21.495 2.475 ;
        RECT 18.155 0.945 18.435 1.405 ;
        RECT 19.450 0.945 19.835 1.515 ;
        RECT 20.540 1.405 21.495 1.575 ;
        RECT 21.665 2.305 22.065 3.155 ;
        RECT 22.255 2.695 22.535 3.155 ;
        RECT 22.255 2.475 23.380 2.695 ;
        RECT 21.665 1.745 22.760 2.305 ;
        RECT 22.930 2.015 23.380 2.475 ;
        RECT 23.550 2.300 23.935 3.155 ;
        RECT 24.640 2.695 24.925 3.155 ;
        RECT 24.640 2.475 25.595 2.695 ;
        RECT 24.525 2.300 25.215 2.305 ;
        RECT 23.550 2.185 25.215 2.300 ;
        RECT 20.540 0.945 20.825 1.405 ;
        RECT 21.665 0.945 22.065 1.745 ;
        RECT 22.930 1.685 23.485 2.015 ;
        RECT 23.655 1.750 25.215 2.185 ;
        RECT 22.930 1.575 23.380 1.685 ;
        RECT 22.255 1.405 23.380 1.575 ;
        RECT 23.655 1.515 23.935 1.750 ;
        RECT 24.525 1.745 25.215 1.750 ;
        RECT 25.385 1.575 25.595 2.475 ;
        RECT 22.255 0.945 22.535 1.405 ;
        RECT 23.550 0.945 23.935 1.515 ;
        RECT 24.640 1.405 25.595 1.575 ;
        RECT 25.765 2.305 26.165 3.155 ;
        RECT 26.355 2.695 26.635 3.155 ;
        RECT 26.355 2.475 27.480 2.695 ;
        RECT 25.765 1.745 26.860 2.305 ;
        RECT 27.030 2.015 27.480 2.475 ;
        RECT 27.650 2.185 28.035 3.155 ;
        RECT 24.640 0.945 24.925 1.405 ;
        RECT 25.765 0.945 26.165 1.745 ;
        RECT 27.030 1.685 27.585 2.015 ;
        RECT 27.030 1.575 27.480 1.685 ;
        RECT 26.355 1.405 27.480 1.575 ;
        RECT 27.755 1.600 28.035 2.185 ;
        RECT 27.755 1.515 29.450 1.600 ;
        RECT 26.355 0.945 26.635 1.405 ;
        RECT 27.650 1.250 29.450 1.515 ;
        RECT 27.650 0.945 28.035 1.250 ;
        RECT 29.100 0.250 29.450 1.250 ;
        RECT 18.500 -0.100 29.450 0.250 ;
        RECT 3.815 -1.605 3.985 -0.845 ;
        RECT 3.815 -1.775 4.530 -1.605 ;
        RECT 4.700 -1.750 4.955 -0.845 ;
        RECT 7.615 -1.345 7.785 -0.845 ;
        RECT 7.615 -1.515 8.280 -1.345 ;
        RECT 4.360 -1.985 4.530 -1.775 ;
        RECT 4.360 -2.315 4.615 -1.985 ;
        RECT 4.360 -2.505 4.530 -2.315 ;
        RECT 4.785 -2.480 4.955 -1.750 ;
        RECT 3.815 -2.675 4.530 -2.505 ;
        RECT 3.815 -3.055 3.985 -2.675 ;
        RECT 4.700 -3.055 4.955 -2.480 ;
        RECT 8.050 -2.505 8.280 -1.515 ;
        RECT 7.615 -2.675 8.280 -2.505 ;
        RECT 7.615 -2.965 7.785 -2.675 ;
        RECT 8.455 -2.965 8.640 -0.845 ;
        RECT 9.315 -1.270 9.565 -0.845 ;
        RECT 9.775 -1.120 10.880 -0.950 ;
        RECT 9.260 -1.400 9.565 -1.270 ;
        RECT 8.810 -2.595 9.090 -1.645 ;
        RECT 9.260 -2.505 9.430 -1.400 ;
        RECT 9.600 -2.185 9.840 -1.590 ;
        RECT 10.010 -1.655 10.540 -1.290 ;
        RECT 10.010 -2.355 10.180 -1.655 ;
        RECT 10.710 -1.735 10.880 -1.120 ;
        RECT 11.390 -1.175 11.640 -0.845 ;
        RECT 11.865 -1.145 12.750 -0.975 ;
        RECT 10.710 -1.825 11.220 -1.735 ;
        RECT 9.260 -2.635 9.485 -2.505 ;
        RECT 9.655 -2.575 10.180 -2.355 ;
        RECT 10.350 -1.995 11.220 -1.825 ;
        RECT 9.315 -2.775 9.485 -2.635 ;
        RECT 10.350 -2.775 10.520 -1.995 ;
        RECT 11.050 -2.065 11.220 -1.995 ;
        RECT 10.730 -2.245 10.930 -2.215 ;
        RECT 11.390 -2.245 11.560 -1.175 ;
        RECT 11.730 -2.065 11.920 -1.345 ;
        RECT 10.730 -2.545 11.560 -2.245 ;
        RECT 12.090 -2.275 12.410 -1.315 ;
        RECT 9.315 -2.945 9.650 -2.775 ;
        RECT 9.845 -2.945 10.520 -2.775 ;
        RECT 11.390 -2.775 11.560 -2.545 ;
        RECT 11.945 -2.605 12.410 -2.275 ;
        RECT 12.580 -1.985 12.750 -1.145 ;
        RECT 13.475 -1.405 13.815 -0.845 ;
        RECT 12.920 -1.780 13.815 -1.405 ;
        RECT 13.625 -1.985 13.815 -1.780 ;
        RECT 17.225 -1.825 17.555 -0.845 ;
        RECT 12.580 -2.315 13.455 -1.985 ;
        RECT 13.625 -2.315 14.375 -1.985 ;
        RECT 12.580 -2.775 12.750 -2.315 ;
        RECT 13.625 -2.485 13.825 -2.315 ;
        RECT 11.390 -2.945 11.795 -2.775 ;
        RECT 11.965 -2.945 12.750 -2.775 ;
        RECT 13.495 -3.010 13.825 -2.485 ;
        RECT 17.290 -2.425 17.460 -1.825 ;
        RECT 17.630 -2.000 17.965 -1.985 ;
        RECT 18.500 -2.000 18.850 -0.100 ;
        RECT 17.630 -2.235 18.850 -2.000 ;
        RECT 19.445 -2.235 19.775 -1.985 ;
        RECT 17.950 -2.250 18.850 -2.235 ;
        RECT 17.290 -3.055 17.985 -2.425 ;
      LAYER met1 ;
        RECT 4.670 -1.860 4.970 -1.010 ;
        RECT 8.010 -1.370 8.300 -1.325 ;
        RECT 10.110 -1.370 10.400 -1.325 ;
        RECT 11.680 -1.370 11.970 -1.325 ;
        RECT 8.010 -1.510 11.970 -1.370 ;
        RECT 8.010 -1.555 8.300 -1.510 ;
        RECT 10.110 -1.555 10.400 -1.510 ;
        RECT 11.680 -1.555 11.970 -1.510 ;
        RECT 4.680 -1.960 4.970 -1.860 ;
        RECT 8.405 -1.710 8.695 -1.665 ;
        RECT 9.595 -1.710 9.885 -1.665 ;
        RECT 12.115 -1.710 12.405 -1.665 ;
        RECT 8.405 -1.850 12.405 -1.710 ;
        RECT 8.405 -1.895 8.695 -1.850 ;
        RECT 9.595 -1.895 9.885 -1.850 ;
        RECT 12.115 -1.895 12.405 -1.850 ;
        RECT 4.680 -2.260 6.560 -1.960 ;
        RECT 6.330 -2.550 6.560 -2.260 ;
        RECT 8.790 -2.550 9.070 -2.260 ;
        RECT 19.050 -2.300 19.800 -1.950 ;
        RECT 19.050 -2.400 19.350 -2.300 ;
        RECT 6.330 -2.850 9.070 -2.550 ;
        RECT 17.300 -2.700 19.350 -2.400 ;
  END
END qz
MACRO vco
  CLASS BLOCK ;
  FOREIGN vco ;
  ORIGIN 0.000 0.000 ;
  SIZE 99.650 BY 36.650 ;
  PIN VCCD
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.841500 ;
    PORT
      LAYER nwell ;
        RECT 25.450 14.500 28.850 16.100 ;
        RECT 25.450 14.495 28.130 14.500 ;
      LAYER li1 ;
        RECT 25.640 15.825 27.940 15.995 ;
        RECT 26.155 15.425 27.090 15.825 ;
        RECT 27.615 14.850 27.855 15.145 ;
        RECT 28.200 15.050 28.600 15.550 ;
        RECT 27.615 14.350 28.050 14.850 ;
        RECT 27.615 14.165 27.855 14.350 ;
      LAYER met1 ;
        RECT 25.550 16.850 29.750 17.350 ;
        RECT 25.650 16.150 26.150 16.850 ;
        RECT 25.640 15.670 27.940 16.150 ;
        RECT 28.200 15.050 28.600 16.850 ;
        RECT 27.450 14.650 28.050 14.950 ;
        RECT 29.250 14.650 29.750 16.850 ;
        RECT 27.450 14.350 29.750 14.650 ;
    END
  END VCCD
  PIN ENB
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 25.725 14.850 26.185 14.915 ;
        RECT 24.950 14.550 26.185 14.850 ;
        RECT 25.725 14.185 26.185 14.550 ;
    END
  END ENB
  PIN p[4]
    ANTENNAGATEAREA 98.549995 ;
    ANTENNADIFFAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 5.100 28.000 6.300 28.650 ;
        RECT 8.800 28.000 10.000 28.650 ;
        RECT 42.700 2.800 43.100 12.850 ;
        RECT 57.650 9.700 58.050 12.850 ;
        RECT 54.700 9.200 58.050 9.700 ;
        RECT 49.850 8.600 51.050 8.650 ;
        RECT 54.700 8.600 55.200 9.200 ;
        RECT 49.850 8.100 55.200 8.600 ;
        RECT 49.850 8.000 51.050 8.100 ;
        RECT 57.650 2.800 58.050 9.200 ;
      LAYER met1 ;
        RECT 0.000 31.750 7.000 32.250 ;
        RECT 0.000 4.900 0.500 31.750 ;
        RECT 6.500 28.650 7.000 31.750 ;
        RECT 5.100 28.000 10.000 28.650 ;
        RECT 49.850 8.000 51.050 8.650 ;
        RECT 42.700 4.900 43.100 5.300 ;
        RECT 50.200 4.900 50.700 8.000 ;
        RECT 57.650 4.900 58.050 5.300 ;
        RECT 0.000 4.400 58.050 4.900 ;
        RECT 42.700 3.900 43.100 4.400 ;
        RECT 57.650 3.900 58.050 4.400 ;
    END
  END p[4]
  PIN Anlg_in
    PORT
      LAYER li1 ;
        RECT 20.830 19.400 21.000 19.480 ;
        RECT 20.830 19.080 22.815 19.400 ;
        RECT 20.830 19.000 21.000 19.080 ;
      LAYER met1 ;
        RECT 20.450 19.430 20.850 19.500 ;
        RECT 20.450 19.050 22.875 19.430 ;
        RECT 20.450 18.950 20.850 19.050 ;
    END
  END Anlg_in
  PIN VCCA
    ANTENNADIFFAREA 4.000000 ;
    PORT
      LAYER nwell ;
        RECT 3.000 28.450 93.000 34.250 ;
        RECT 33.000 2.400 93.000 8.200 ;
      LAYER li1 ;
        RECT 3.200 33.400 3.600 33.900 ;
        RECT 12.700 33.400 13.100 33.900 ;
        RECT 18.150 33.400 18.550 33.900 ;
        RECT 23.600 33.400 24.000 33.900 ;
        RECT 33.200 33.400 33.600 33.900 ;
        RECT 42.700 33.400 43.100 33.900 ;
        RECT 48.150 33.400 48.550 33.900 ;
        RECT 53.600 33.400 54.000 33.900 ;
        RECT 63.200 33.400 63.600 33.900 ;
        RECT 72.700 33.400 73.100 33.900 ;
        RECT 78.150 33.400 78.550 33.900 ;
        RECT 83.600 33.400 84.000 33.900 ;
        RECT 42.000 2.750 42.400 3.250 ;
        RECT 47.450 2.750 47.850 3.250 ;
        RECT 52.900 2.750 53.300 3.250 ;
        RECT 62.400 2.750 62.800 3.250 ;
        RECT 72.000 2.750 72.400 3.250 ;
        RECT 77.450 2.750 77.850 3.250 ;
        RECT 82.900 2.750 83.300 3.250 ;
        RECT 92.400 2.750 92.800 3.250 ;
      LAYER met1 ;
        RECT 3.200 36.150 99.650 36.650 ;
        RECT 3.200 33.400 3.600 36.150 ;
        RECT 12.700 33.400 13.100 36.150 ;
        RECT 18.150 33.400 18.550 36.150 ;
        RECT 23.600 33.400 24.000 36.150 ;
        RECT 33.200 33.400 33.600 36.150 ;
        RECT 42.700 33.400 43.100 36.150 ;
        RECT 48.150 33.400 48.550 36.150 ;
        RECT 53.600 33.400 54.000 36.150 ;
        RECT 63.200 33.400 63.600 36.150 ;
        RECT 72.700 33.400 73.100 36.150 ;
        RECT 78.150 33.400 78.550 36.150 ;
        RECT 83.600 33.400 84.000 36.150 ;
        RECT 42.000 0.500 42.400 3.250 ;
        RECT 47.450 0.500 47.850 3.250 ;
        RECT 52.900 0.500 53.300 3.250 ;
        RECT 62.400 0.500 62.800 3.250 ;
        RECT 72.000 0.500 72.400 3.250 ;
        RECT 77.450 0.500 77.850 3.250 ;
        RECT 82.900 0.500 83.300 3.250 ;
        RECT 92.400 0.500 92.800 3.250 ;
        RECT 97.050 0.500 97.550 36.150 ;
        RECT 42.000 0.000 97.550 0.500 ;
    END
  END VCCA
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 3.900 34.750 99.650 35.150 ;
        RECT 3.900 28.850 4.300 34.750 ;
        RECT 12.000 28.850 12.400 34.750 ;
        RECT 13.400 28.850 13.800 34.750 ;
        RECT 18.850 28.850 19.250 34.750 ;
        RECT 24.300 28.850 24.700 34.750 ;
        RECT 32.400 28.850 32.800 34.750 ;
        RECT 33.900 28.850 34.300 34.750 ;
        RECT 42.000 28.850 42.400 34.750 ;
        RECT 43.400 28.850 43.800 34.750 ;
        RECT 48.850 28.850 49.250 34.750 ;
        RECT 54.300 28.850 54.700 34.750 ;
        RECT 62.400 28.850 62.800 34.750 ;
        RECT 63.900 28.850 64.300 34.750 ;
        RECT 72.000 28.850 72.400 34.750 ;
        RECT 73.400 28.850 73.800 34.750 ;
        RECT 78.850 28.850 79.250 34.750 ;
        RECT 84.300 28.850 84.700 34.750 ;
        RECT 92.400 28.850 92.800 34.750 ;
        RECT 33.200 1.900 33.600 7.800 ;
        RECT 41.300 1.900 41.700 7.800 ;
        RECT 46.750 1.900 47.150 7.800 ;
        RECT 52.200 1.900 52.600 7.800 ;
        RECT 53.600 1.900 54.000 7.800 ;
        RECT 61.700 1.900 62.100 7.800 ;
        RECT 63.200 1.900 63.600 7.800 ;
        RECT 71.300 1.900 71.700 7.800 ;
        RECT 76.750 1.900 77.150 7.800 ;
        RECT 82.200 1.900 82.600 7.800 ;
        RECT 83.600 1.900 84.000 7.800 ;
        RECT 91.700 1.900 92.100 7.800 ;
        RECT 98.550 1.900 99.050 34.750 ;
        RECT 33.200 1.500 99.050 1.900 ;
    END
  END VPWR
  PIN GND
    ANTENNADIFFAREA 4.394000 ;
    PORT
      LAYER pwell ;
        RECT 3.000 23.400 93.000 28.200 ;
        RECT 26.130 14.200 27.935 14.205 ;
        RECT 26.130 13.975 28.850 14.200 ;
        RECT 25.645 13.300 28.850 13.975 ;
        RECT 25.645 13.295 27.935 13.300 ;
        RECT 25.790 13.105 25.960 13.295 ;
        RECT 33.000 8.450 93.000 13.250 ;
      LAYER li1 ;
        RECT 3.200 23.750 3.600 24.250 ;
        RECT 12.700 23.750 13.100 24.250 ;
        RECT 18.150 23.750 18.550 24.250 ;
        RECT 23.600 23.750 24.000 24.250 ;
        RECT 33.200 23.750 33.600 24.250 ;
        RECT 42.700 23.750 43.100 24.250 ;
        RECT 48.150 23.750 48.550 24.250 ;
        RECT 53.600 23.750 54.000 24.250 ;
        RECT 63.200 23.750 63.600 24.250 ;
        RECT 72.700 23.750 73.100 24.250 ;
        RECT 78.150 23.750 78.550 24.250 ;
        RECT 83.600 23.750 84.000 24.250 ;
        RECT 41.100 17.850 41.270 17.930 ;
        RECT 39.285 17.530 41.270 17.850 ;
        RECT 41.100 17.450 41.270 17.530 ;
        RECT 26.155 13.275 27.090 13.675 ;
        RECT 28.200 13.550 28.600 14.050 ;
        RECT 25.640 13.105 27.940 13.275 ;
        RECT 42.000 12.400 42.400 12.900 ;
        RECT 47.450 12.400 47.850 12.900 ;
        RECT 52.900 12.400 53.300 12.900 ;
        RECT 62.400 12.400 62.800 12.900 ;
        RECT 72.000 12.400 72.400 12.900 ;
        RECT 77.450 12.400 77.850 12.900 ;
        RECT 82.900 12.400 83.300 12.900 ;
        RECT 92.400 12.400 92.800 12.900 ;
      LAYER met1 ;
        RECT 3.200 21.500 3.600 24.250 ;
        RECT 12.700 21.500 13.100 24.250 ;
        RECT 18.150 21.500 18.550 24.250 ;
        RECT 23.600 21.500 24.000 24.250 ;
        RECT 33.200 21.500 33.600 24.250 ;
        RECT 42.700 21.500 43.100 24.250 ;
        RECT 48.150 21.500 48.550 24.250 ;
        RECT 53.600 21.500 54.000 24.250 ;
        RECT 63.200 21.500 63.600 24.250 ;
        RECT 72.700 21.500 73.100 24.250 ;
        RECT 78.150 21.500 78.550 24.250 ;
        RECT 83.600 21.500 84.000 24.250 ;
        RECT 3.200 21.000 84.000 21.500 ;
        RECT 28.200 13.900 28.600 14.050 ;
        RECT 31.150 13.900 31.650 21.000 ;
        RECT 42.000 17.950 42.500 21.000 ;
        RECT 41.150 17.880 42.500 17.950 ;
        RECT 39.225 17.500 42.500 17.880 ;
        RECT 41.150 17.400 42.500 17.500 ;
        RECT 28.200 13.600 31.650 13.900 ;
        RECT 28.200 13.550 28.600 13.600 ;
        RECT 25.640 13.250 27.940 13.430 ;
        RECT 31.150 13.250 31.650 13.600 ;
        RECT 25.640 12.950 31.650 13.250 ;
        RECT 42.000 15.650 42.500 17.400 ;
        RECT 83.500 15.650 84.000 21.000 ;
        RECT 42.000 15.150 92.800 15.650 ;
        RECT 42.000 12.400 42.400 15.150 ;
        RECT 47.450 12.400 47.850 15.150 ;
        RECT 52.900 12.400 53.300 15.150 ;
        RECT 62.400 12.400 62.800 15.150 ;
        RECT 72.000 12.400 72.400 15.150 ;
        RECT 77.450 12.400 77.850 15.150 ;
        RECT 82.900 12.400 83.300 15.150 ;
        RECT 92.400 12.400 92.800 15.150 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 3.900 22.900 4.300 27.800 ;
        RECT 7.950 27.450 8.350 33.850 ;
        RECT 14.950 28.550 16.150 28.650 ;
        RECT 10.800 28.050 16.150 28.550 ;
        RECT 10.800 27.450 11.300 28.050 ;
        RECT 14.950 28.000 16.150 28.050 ;
        RECT 17.450 28.600 17.850 33.850 ;
        RECT 19.800 28.600 21.000 28.650 ;
        RECT 17.450 28.100 21.000 28.600 ;
        RECT 7.950 26.950 11.300 27.450 ;
        RECT 7.950 23.800 8.350 26.950 ;
        RECT 12.000 22.900 12.400 27.800 ;
        RECT 13.400 22.900 13.800 27.800 ;
        RECT 17.450 23.800 17.850 28.100 ;
        RECT 19.800 28.000 21.000 28.100 ;
        RECT 18.850 22.900 19.250 27.800 ;
        RECT 22.900 23.800 23.300 33.850 ;
        RECT 25.500 28.000 26.700 28.650 ;
        RECT 24.300 22.900 24.700 27.800 ;
        RECT 28.350 23.800 28.750 33.850 ;
        RECT 29.200 28.000 30.400 28.650 ;
        RECT 35.100 28.000 36.300 28.650 ;
        RECT 32.400 22.900 32.800 27.800 ;
        RECT 33.900 22.900 34.300 27.800 ;
        RECT 37.950 27.450 38.350 33.850 ;
        RECT 38.800 28.000 40.000 28.650 ;
        RECT 44.950 28.550 46.150 28.650 ;
        RECT 40.800 28.050 46.150 28.550 ;
        RECT 40.800 27.450 41.300 28.050 ;
        RECT 44.950 28.000 46.150 28.050 ;
        RECT 47.450 28.600 47.850 33.850 ;
        RECT 49.800 28.600 51.000 28.650 ;
        RECT 47.450 28.100 51.000 28.600 ;
        RECT 37.950 26.950 41.300 27.450 ;
        RECT 37.950 23.800 38.350 26.950 ;
        RECT 42.000 22.900 42.400 27.800 ;
        RECT 43.400 22.900 43.800 27.800 ;
        RECT 47.450 23.800 47.850 28.100 ;
        RECT 49.800 28.000 51.000 28.100 ;
        RECT 48.850 22.900 49.250 27.800 ;
        RECT 52.900 23.800 53.300 33.850 ;
        RECT 55.500 28.000 56.700 28.650 ;
        RECT 54.300 22.900 54.700 27.800 ;
        RECT 58.350 23.800 58.750 33.850 ;
        RECT 59.200 28.000 60.400 28.650 ;
        RECT 65.100 28.000 66.300 28.650 ;
        RECT 62.400 22.900 62.800 27.800 ;
        RECT 63.900 22.900 64.300 27.800 ;
        RECT 67.950 27.450 68.350 33.850 ;
        RECT 68.800 28.000 70.000 28.650 ;
        RECT 74.950 28.550 76.150 28.650 ;
        RECT 70.800 28.050 76.150 28.550 ;
        RECT 70.800 27.450 71.300 28.050 ;
        RECT 74.950 28.000 76.150 28.050 ;
        RECT 77.450 28.600 77.850 33.850 ;
        RECT 79.800 28.600 81.000 28.650 ;
        RECT 77.450 28.100 81.000 28.600 ;
        RECT 67.950 26.950 71.300 27.450 ;
        RECT 67.950 23.800 68.350 26.950 ;
        RECT 72.000 22.900 72.400 27.800 ;
        RECT 73.400 22.900 73.800 27.800 ;
        RECT 77.450 23.800 77.850 28.100 ;
        RECT 79.800 28.000 81.000 28.100 ;
        RECT 78.850 22.900 79.250 27.800 ;
        RECT 82.900 23.800 83.300 33.850 ;
        RECT 85.500 28.000 86.700 28.650 ;
        RECT 84.300 22.900 84.700 27.800 ;
        RECT 88.350 23.800 88.750 33.850 ;
        RECT 89.200 28.000 90.400 28.650 ;
        RECT 92.400 22.900 92.800 27.800 ;
        RECT 3.900 22.500 92.800 22.900 ;
        RECT 26.950 19.480 27.350 19.500 ;
        RECT 26.800 19.450 27.350 19.480 ;
        RECT 33.950 19.450 34.450 22.500 ;
        RECT 26.800 19.400 34.450 19.450 ;
        RECT 24.985 19.080 34.450 19.400 ;
        RECT 26.800 19.050 34.450 19.080 ;
        RECT 26.800 19.000 27.350 19.050 ;
        RECT 33.950 18.000 34.450 19.050 ;
        RECT 33.950 17.930 35.200 18.000 ;
        RECT 33.950 17.850 35.300 17.930 ;
        RECT 33.950 17.530 37.115 17.850 ;
        RECT 33.950 17.450 35.300 17.530 ;
        RECT 33.950 17.400 35.200 17.450 ;
        RECT 25.725 15.255 25.985 15.655 ;
        RECT 27.260 15.315 27.855 15.655 ;
        RECT 25.725 15.085 27.090 15.255 ;
        RECT 26.355 14.015 27.090 15.085 ;
        RECT 25.725 13.845 27.090 14.015 ;
        RECT 27.260 13.995 27.435 15.315 ;
        RECT 33.950 14.150 34.450 17.400 ;
        RECT 91.600 14.150 92.100 22.500 ;
        RECT 25.725 13.445 25.985 13.845 ;
        RECT 27.260 13.445 27.855 13.995 ;
        RECT 33.200 13.750 92.100 14.150 ;
        RECT 33.200 8.850 33.600 13.750 ;
        RECT 35.600 8.000 36.800 8.650 ;
        RECT 37.250 2.800 37.650 12.850 ;
        RECT 41.300 8.850 41.700 13.750 ;
        RECT 46.750 8.850 47.150 13.750 ;
        RECT 39.300 8.000 40.500 8.650 ;
        RECT 45.000 8.550 46.200 8.650 ;
        RECT 48.150 8.550 48.550 12.850 ;
        RECT 52.200 8.850 52.600 13.750 ;
        RECT 53.600 8.850 54.000 13.750 ;
        RECT 61.700 8.850 62.100 13.750 ;
        RECT 63.200 8.850 63.600 13.750 ;
        RECT 45.000 8.050 48.550 8.550 ;
        RECT 45.000 8.000 46.200 8.050 ;
        RECT 48.150 2.800 48.550 8.050 ;
        RECT 56.000 8.000 57.200 8.650 ;
        RECT 59.700 8.000 60.900 8.650 ;
        RECT 65.600 8.000 66.800 8.650 ;
        RECT 67.250 2.800 67.650 12.850 ;
        RECT 71.300 8.850 71.700 13.750 ;
        RECT 69.300 8.000 70.500 8.650 ;
        RECT 72.700 2.800 73.100 12.850 ;
        RECT 76.750 8.850 77.150 13.750 ;
        RECT 75.000 8.550 76.200 8.650 ;
        RECT 78.150 8.550 78.550 12.850 ;
        RECT 82.200 8.850 82.600 13.750 ;
        RECT 83.600 8.850 84.000 13.750 ;
        RECT 87.650 9.700 88.050 12.850 ;
        RECT 84.700 9.200 88.050 9.700 ;
        RECT 75.000 8.050 78.550 8.550 ;
        RECT 75.000 8.000 76.200 8.050 ;
        RECT 78.150 2.800 78.550 8.050 ;
        RECT 79.850 8.600 81.050 8.650 ;
        RECT 84.700 8.600 85.200 9.200 ;
        RECT 79.850 8.100 85.200 8.600 ;
        RECT 79.850 8.000 81.050 8.100 ;
        RECT 86.000 8.000 87.200 8.650 ;
        RECT 87.650 2.800 88.050 9.200 ;
        RECT 91.700 8.850 92.100 13.750 ;
        RECT 89.700 8.000 90.900 8.650 ;
      LAYER met1 ;
        RECT 7.950 32.250 8.350 32.750 ;
        RECT 22.900 32.250 23.300 32.750 ;
        RECT 37.950 32.250 38.350 32.750 ;
        RECT 52.900 32.250 53.300 32.750 ;
        RECT 67.950 32.250 68.350 32.750 ;
        RECT 82.900 32.250 83.300 32.750 ;
        RECT 7.950 31.750 37.000 32.250 ;
        RECT 7.950 31.350 8.350 31.750 ;
        RECT 15.300 28.650 15.800 31.750 ;
        RECT 22.900 31.350 23.300 31.750 ;
        RECT 17.450 30.700 17.850 31.050 ;
        RECT 28.350 30.700 28.750 31.050 ;
        RECT 17.450 30.200 28.750 30.700 ;
        RECT 17.450 29.850 17.850 30.200 ;
        RECT 20.150 28.650 20.650 30.200 ;
        RECT 28.350 29.850 28.750 30.200 ;
        RECT 36.500 28.650 37.000 31.750 ;
        RECT 37.950 31.750 67.000 32.250 ;
        RECT 37.950 31.350 38.350 31.750 ;
        RECT 45.300 28.650 45.800 31.750 ;
        RECT 52.900 31.350 53.300 31.750 ;
        RECT 47.450 30.700 47.850 31.050 ;
        RECT 58.350 30.700 58.750 31.050 ;
        RECT 47.450 30.200 58.750 30.700 ;
        RECT 47.450 29.850 47.850 30.200 ;
        RECT 50.150 28.650 50.650 30.200 ;
        RECT 58.350 29.850 58.750 30.200 ;
        RECT 66.500 28.650 67.000 31.750 ;
        RECT 67.950 31.750 96.000 32.250 ;
        RECT 67.950 31.350 68.350 31.750 ;
        RECT 75.300 28.650 75.800 31.750 ;
        RECT 82.900 31.350 83.300 31.750 ;
        RECT 77.450 30.700 77.850 31.050 ;
        RECT 88.350 30.700 88.750 31.050 ;
        RECT 77.450 30.200 88.750 30.700 ;
        RECT 77.450 29.850 77.850 30.200 ;
        RECT 80.150 28.650 80.650 30.200 ;
        RECT 88.350 29.850 88.750 30.200 ;
        RECT 14.950 28.000 16.150 28.650 ;
        RECT 19.800 28.000 21.000 28.650 ;
        RECT 25.500 28.550 30.400 28.650 ;
        RECT 24.650 28.050 30.400 28.550 ;
        RECT 24.650 25.900 25.150 28.050 ;
        RECT 25.500 28.000 30.400 28.050 ;
        RECT 35.100 28.000 40.000 28.650 ;
        RECT 44.950 28.000 46.150 28.650 ;
        RECT 49.800 28.000 51.000 28.650 ;
        RECT 55.500 28.550 60.400 28.650 ;
        RECT 54.650 28.050 60.400 28.550 ;
        RECT 1.500 25.400 25.150 25.900 ;
        RECT 28.350 25.900 28.750 26.200 ;
        RECT 54.650 25.900 55.150 28.050 ;
        RECT 55.500 28.000 60.400 28.050 ;
        RECT 65.100 28.000 70.000 28.650 ;
        RECT 74.950 28.000 76.150 28.650 ;
        RECT 79.800 28.000 81.000 28.650 ;
        RECT 85.500 28.550 90.400 28.650 ;
        RECT 84.650 28.050 90.400 28.550 ;
        RECT 28.350 25.400 55.150 25.900 ;
        RECT 58.350 25.900 58.750 26.200 ;
        RECT 84.650 25.900 85.150 28.050 ;
        RECT 85.500 28.000 90.400 28.050 ;
        RECT 58.350 25.400 85.150 25.900 ;
        RECT 88.350 25.900 88.750 26.200 ;
        RECT 88.350 25.400 94.500 25.900 ;
        RECT 1.500 11.250 2.000 25.400 ;
        RECT 28.350 25.000 28.750 25.400 ;
        RECT 58.350 25.000 58.750 25.400 ;
        RECT 88.350 25.000 88.750 25.400 ;
        RECT 24.925 19.050 27.030 19.430 ;
        RECT 35.070 17.500 37.175 17.880 ;
        RECT 27.400 14.000 27.850 14.100 ;
        RECT 24.450 13.700 27.850 14.000 ;
        RECT 24.450 11.250 24.950 13.700 ;
        RECT 27.400 13.650 27.850 13.700 ;
        RECT 37.250 11.250 37.650 11.650 ;
        RECT 67.250 11.250 67.650 11.650 ;
        RECT 94.000 11.250 94.500 25.400 ;
        RECT 1.500 10.750 37.650 11.250 ;
        RECT 37.250 10.450 37.650 10.750 ;
        RECT 40.850 10.750 67.650 11.250 ;
        RECT 35.600 8.600 40.500 8.650 ;
        RECT 40.850 8.600 41.350 10.750 ;
        RECT 67.250 10.450 67.650 10.750 ;
        RECT 70.850 10.750 94.500 11.250 ;
        RECT 35.600 8.100 41.350 8.600 ;
        RECT 35.600 8.000 40.500 8.100 ;
        RECT 45.000 8.000 46.200 8.650 ;
        RECT 56.000 8.000 60.900 8.650 ;
        RECT 65.600 8.600 70.500 8.650 ;
        RECT 70.850 8.600 71.350 10.750 ;
        RECT 65.600 8.100 71.350 8.600 ;
        RECT 65.600 8.000 70.500 8.100 ;
        RECT 75.000 8.000 76.200 8.650 ;
        RECT 79.850 8.000 81.050 8.650 ;
        RECT 86.000 8.000 90.900 8.650 ;
        RECT 37.250 6.450 37.650 6.800 ;
        RECT 45.350 6.450 45.850 8.000 ;
        RECT 48.150 6.450 48.550 6.800 ;
        RECT 37.250 5.950 48.550 6.450 ;
        RECT 37.250 5.600 37.650 5.950 ;
        RECT 48.150 5.600 48.550 5.950 ;
        RECT 59.000 4.900 59.500 8.000 ;
        RECT 67.250 6.450 67.650 6.800 ;
        RECT 75.350 6.450 75.850 8.000 ;
        RECT 78.150 6.450 78.550 6.800 ;
        RECT 67.250 5.950 78.550 6.450 ;
        RECT 67.250 5.600 67.650 5.950 ;
        RECT 78.150 5.600 78.550 5.950 ;
        RECT 72.700 4.900 73.100 5.300 ;
        RECT 80.200 4.900 80.700 8.000 ;
        RECT 87.650 4.900 88.050 5.300 ;
        RECT 59.000 4.400 88.050 4.900 ;
        RECT 89.000 4.900 89.500 8.000 ;
        RECT 95.500 4.900 96.000 31.750 ;
        RECT 89.000 4.400 96.000 4.900 ;
        RECT 72.700 3.900 73.100 4.400 ;
        RECT 87.650 3.900 88.050 4.400 ;
  END
END vco
MACRO system
  CLASS BLOCK ;
  FOREIGN system ;
  ORIGIN 26.425 62.950 ;
  SIZE 134.975 BY 103.000 ;
  PIN Dout
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 90.625 -12.885 90.955 -12.040 ;
        RECT 90.625 -12.965 91.015 -12.885 ;
        RECT 90.800 -13.015 91.015 -12.965 ;
        RECT 90.845 -13.150 91.015 -13.015 ;
        RECT 93.085 -13.150 93.420 -13.135 ;
        RECT 90.845 -13.400 93.420 -13.150 ;
        RECT 90.845 -13.595 91.015 -13.400 ;
        RECT 90.790 -13.635 91.015 -13.595 ;
        RECT 90.635 -13.720 91.015 -13.635 ;
        RECT 90.635 -14.155 90.965 -13.720 ;
        RECT 92.000 -16.000 92.350 -13.400 ;
        RECT 93.085 -13.405 93.420 -13.400 ;
    END
  END Dout
  PIN CLK
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER li1 ;
        RECT 78.500 -9.300 78.850 -5.350 ;
        RECT 80.025 -9.405 80.715 -8.845 ;
        RECT 83.830 -13.485 84.180 -12.835 ;
      LAYER met1 ;
        RECT 80.030 -8.950 80.730 -8.830 ;
        RECT 78.500 -9.300 80.730 -8.950 ;
        RECT 78.500 -10.950 78.850 -9.300 ;
        RECT 80.030 -9.400 80.730 -9.300 ;
        RECT 78.500 -11.300 83.350 -10.950 ;
        RECT 83.000 -12.800 83.350 -11.300 ;
        RECT 83.000 -12.840 84.150 -12.800 ;
        RECT 83.000 -13.150 84.160 -12.840 ;
        RECT 83.810 -13.490 84.160 -13.150 ;
    END
  END CLK
  PIN Anlg_in
    PORT
      LAYER li1 ;
        RECT -13.800 22.880 10.750 22.900 ;
        RECT -13.800 22.800 10.900 22.880 ;
        RECT -13.800 22.480 12.715 22.800 ;
        RECT -13.800 22.400 10.900 22.480 ;
        RECT -13.800 22.350 10.750 22.400 ;
      LAYER met1 ;
        RECT 10.350 22.830 10.750 22.900 ;
        RECT 10.350 22.450 12.775 22.830 ;
        RECT 10.350 22.350 10.750 22.450 ;
    END
  END Anlg_in
  PIN VCCD
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 33.665051 ;
    PORT
      LAYER nwell ;
        RECT 15.350 17.900 18.750 19.500 ;
        RECT 15.350 17.895 18.030 17.900 ;
        RECT 79.950 -7.550 104.650 -7.500 ;
        RECT 79.750 -9.200 104.650 -7.550 ;
        RECT 80.900 -11.550 97.250 -11.500 ;
        RECT -16.000 -14.280 1.750 -12.580 ;
        RECT 79.750 -13.200 97.250 -11.550 ;
        RECT 28.500 -16.750 32.030 -15.150 ;
        RECT 29.350 -16.755 32.030 -16.750 ;
        RECT -15.950 -17.840 -15.050 -17.780 ;
        RECT -15.950 -19.445 -13.490 -17.840 ;
        RECT -3.650 -18.310 -2.650 -18.280 ;
        RECT -15.950 -19.480 -15.100 -19.445 ;
        RECT -7.240 -19.915 -0.440 -18.310 ;
        RECT -3.650 -19.930 -2.650 -19.915 ;
        RECT -12.650 -24.495 -11.800 -24.480 ;
        RECT -1.900 -24.495 -0.100 -24.480 ;
        RECT -14.390 -26.100 1.890 -24.495 ;
        RECT -12.650 -26.130 -11.800 -26.100 ;
        RECT -1.900 -26.130 0.050 -26.100 ;
        RECT 46.950 -29.750 49.800 -28.150 ;
        RECT 46.950 -29.755 49.170 -29.750 ;
        RECT 52.650 -30.850 54.800 -30.800 ;
        RECT 52.650 -32.450 67.040 -30.850 ;
        RECT 54.700 -32.455 67.040 -32.450 ;
        RECT 57.300 -32.500 59.400 -32.455 ;
        RECT 51.650 -36.650 69.400 -35.050 ;
        RECT 77.350 -36.330 95.100 -34.630 ;
        RECT 52.500 -36.655 69.400 -36.650 ;
        RECT 55.600 -36.700 57.950 -36.655 ;
        RECT 67.900 -36.700 69.400 -36.655 ;
        RECT 77.400 -39.890 78.300 -39.830 ;
        RECT 77.400 -41.495 79.860 -39.890 ;
        RECT 89.700 -40.360 90.700 -40.330 ;
        RECT 77.400 -41.530 78.250 -41.495 ;
        RECT 19.645 -43.950 21.250 -41.800 ;
        RECT 86.110 -41.965 92.910 -40.360 ;
        RECT 89.700 -41.980 90.700 -41.965 ;
        RECT 19.600 -45.100 21.250 -43.950 ;
        RECT 52.650 -42.550 54.800 -42.500 ;
        RECT 52.650 -44.150 67.040 -42.550 ;
        RECT 54.700 -44.155 67.040 -44.150 ;
        RECT 57.300 -44.200 59.400 -44.155 ;
        RECT 19.645 -46.860 21.250 -45.100 ;
        RECT 80.700 -46.545 81.550 -46.530 ;
        RECT 91.450 -46.545 93.250 -46.530 ;
        RECT 51.650 -48.350 69.400 -46.750 ;
        RECT 78.960 -48.150 95.240 -46.545 ;
        RECT 80.700 -48.180 81.550 -48.150 ;
        RECT 91.450 -48.180 93.400 -48.150 ;
        RECT 52.500 -48.355 69.400 -48.350 ;
        RECT 55.600 -48.400 57.950 -48.355 ;
        RECT 67.900 -48.400 69.400 -48.355 ;
      LAYER li1 ;
        RECT -13.700 20.750 -12.400 21.350 ;
        RECT -13.700 20.250 16.100 20.750 ;
        RECT -13.700 20.050 -12.400 20.250 ;
        RECT 15.540 19.225 17.840 19.395 ;
        RECT 16.055 18.825 16.990 19.225 ;
        RECT 17.515 18.250 17.755 18.545 ;
        RECT 18.100 18.450 18.500 18.950 ;
        RECT 17.515 17.750 17.950 18.250 ;
        RECT 17.515 17.565 17.755 17.750 ;
        RECT 79.950 -7.655 80.350 -7.500 ;
        RECT 79.940 -7.825 83.620 -7.655 ;
        RECT 84.040 -7.825 87.720 -7.655 ;
        RECT 88.140 -7.825 91.820 -7.655 ;
        RECT 92.540 -7.825 96.220 -7.655 ;
        RECT 96.640 -7.825 100.320 -7.655 ;
        RECT 100.740 -7.825 104.420 -7.655 ;
        RECT 80.595 -8.285 80.865 -7.825 ;
        RECT 82.655 -8.285 82.980 -7.825 ;
        RECT 84.695 -8.285 84.965 -7.825 ;
        RECT 86.755 -8.285 87.080 -7.825 ;
        RECT 88.795 -8.285 89.065 -7.825 ;
        RECT 90.855 -8.285 91.180 -7.825 ;
        RECT 92.050 -8.650 92.450 -8.150 ;
        RECT 93.195 -8.285 93.465 -7.825 ;
        RECT 95.255 -8.285 95.580 -7.825 ;
        RECT 97.295 -8.285 97.565 -7.825 ;
        RECT 99.355 -8.285 99.680 -7.825 ;
        RECT 101.395 -8.285 101.665 -7.825 ;
        RECT 103.455 -8.285 103.780 -7.825 ;
        RECT 81.400 -11.655 84.150 -11.500 ;
        RECT 79.940 -11.700 91.100 -11.655 ;
        RECT 79.940 -11.825 81.780 -11.700 ;
        RECT 80.500 -12.585 80.830 -11.825 ;
        RECT 1.450 -12.735 4.000 -12.730 ;
        RECT -15.210 -12.905 -13.370 -12.735 ;
        RECT -11.770 -12.905 -2.110 -12.735 ;
        RECT -0.300 -12.905 4.000 -12.735 ;
        RECT -14.650 -13.665 -14.320 -12.905 ;
        RECT -13.720 -14.055 -13.460 -12.905 ;
        RECT -12.750 -13.680 -12.350 -13.180 ;
        RECT -11.255 -13.405 -10.925 -12.905 ;
        RECT -10.315 -13.405 -9.985 -12.905 ;
        RECT -8.340 -13.285 -7.960 -12.905 ;
        RECT -7.440 -13.285 -7.110 -12.905 ;
        RECT -5.830 -13.285 -5.410 -12.905 ;
        RECT -4.740 -13.595 -4.410 -12.905 ;
        RECT -3.290 -13.705 -3.005 -12.905 ;
        RECT 0.260 -13.665 0.590 -12.905 ;
        RECT 1.190 -13.080 4.000 -12.905 ;
        RECT 81.430 -12.975 81.690 -11.825 ;
        RECT 82.200 -12.650 82.600 -11.700 ;
        RECT 83.740 -11.825 91.100 -11.700 ;
        RECT 92.990 -11.825 94.370 -11.655 ;
        RECT 95.640 -11.825 97.020 -11.655 ;
        RECT 84.255 -12.325 84.585 -11.825 ;
        RECT 85.180 -12.285 85.445 -11.825 ;
        RECT 87.350 -12.625 87.520 -11.825 ;
        RECT 89.230 -12.325 89.545 -11.825 ;
        RECT 90.285 -12.835 90.455 -11.825 ;
        RECT 93.075 -12.965 93.355 -11.825 ;
        RECT 94.025 -12.965 94.285 -11.825 ;
        RECT 95.765 -12.965 95.995 -11.825 ;
        RECT 96.665 -12.965 96.875 -11.825 ;
        RECT 1.190 -14.055 1.450 -13.080 ;
        RECT -13.850 -17.945 -6.700 -17.930 ;
        RECT -15.060 -18.115 -6.700 -17.945 ;
        RECT -15.750 -18.730 -15.350 -18.230 ;
        RECT -14.935 -19.255 -14.705 -18.115 ;
        RECT -14.035 -18.280 -6.700 -18.115 ;
        RECT -14.035 -19.255 -13.825 -18.280 ;
        RECT -7.050 -18.415 -6.700 -18.280 ;
        RECT -7.050 -18.585 -3.830 -18.415 ;
        RECT -2.470 -18.430 -0.630 -18.415 ;
        RECT 3.650 -18.430 4.000 -13.080 ;
        RECT 29.540 -15.425 31.840 -15.255 ;
        RECT 28.900 -16.270 29.200 -15.770 ;
        RECT 30.055 -15.825 30.990 -15.425 ;
        RECT 31.515 -16.750 31.755 -16.105 ;
        RECT 31.515 -17.050 31.900 -16.750 ;
        RECT 31.515 -17.085 31.755 -17.050 ;
        RECT -2.470 -18.585 4.000 -18.430 ;
        RECT -5.995 -19.435 -5.825 -18.585 ;
        RECT -5.155 -19.095 -4.985 -18.585 ;
        RECT -3.300 -19.480 -2.900 -18.980 ;
        RECT -1.910 -19.345 -1.580 -18.585 ;
        RECT -0.980 -18.780 4.000 -18.585 ;
        RECT -0.980 -19.735 -0.720 -18.780 ;
        RECT -14.055 -25.825 -13.845 -24.685 ;
        RECT -13.175 -25.825 -12.945 -24.685 ;
        RECT -12.350 -25.430 -11.950 -24.930 ;
        RECT -10.835 -25.825 -10.550 -25.025 ;
        RECT -9.430 -25.825 -9.100 -25.135 ;
        RECT -8.430 -25.825 -8.010 -25.445 ;
        RECT -6.730 -25.825 -6.400 -25.445 ;
        RECT -5.880 -25.825 -5.500 -25.445 ;
        RECT -3.855 -25.825 -3.525 -25.325 ;
        RECT -2.915 -25.825 -2.585 -25.325 ;
        RECT -0.050 -25.825 0.210 -24.675 ;
        RECT 0.810 -25.825 1.140 -25.065 ;
        RECT 3.650 -25.780 4.000 -18.780 ;
        RECT 1.650 -25.825 4.000 -25.780 ;
        RECT -14.200 -25.995 -12.820 -25.825 ;
        RECT -11.730 -25.995 -2.070 -25.825 ;
        RECT -0.140 -25.995 4.000 -25.825 ;
        RECT 1.650 -26.130 4.000 -25.995 ;
        RECT 52.850 -27.800 55.400 -27.300 ;
        RECT 47.140 -28.425 48.980 -28.255 ;
        RECT 47.700 -29.185 48.030 -28.425 ;
        RECT 48.630 -29.575 48.890 -28.425 ;
        RECT 49.250 -29.500 49.550 -29.000 ;
        RECT 52.850 -31.850 53.350 -27.800 ;
        RECT 54.900 -30.955 55.400 -27.800 ;
        RECT 66.800 -30.955 68.150 -30.800 ;
        RECT 54.890 -31.125 57.190 -30.955 ;
        RECT 59.490 -31.125 68.150 -30.955 ;
        RECT 55.020 -32.265 55.285 -31.125 ;
        RECT 55.955 -31.925 56.125 -31.125 ;
        RECT 56.795 -31.585 57.005 -31.125 ;
        RECT 60.005 -31.625 60.335 -31.125 ;
        RECT 60.930 -31.585 61.195 -31.125 ;
        RECT 63.100 -31.925 63.270 -31.125 ;
        RECT 64.980 -31.625 65.295 -31.125 ;
        RECT 66.035 -32.135 66.205 -31.125 ;
        RECT 66.800 -31.150 68.150 -31.125 ;
        RECT 67.750 -34.900 68.150 -31.150 ;
        RECT 94.800 -34.785 97.350 -34.780 ;
        RECT 78.140 -34.955 79.980 -34.785 ;
        RECT 81.580 -34.955 91.240 -34.785 ;
        RECT 93.050 -34.955 97.350 -34.785 ;
        RECT 55.450 -35.155 57.100 -35.000 ;
        RECT 52.690 -35.325 57.100 -35.155 ;
        RECT 58.090 -35.325 67.750 -35.155 ;
        RECT 51.950 -36.100 52.350 -35.600 ;
        RECT 53.285 -36.125 53.525 -35.325 ;
        RECT 54.045 -36.125 54.375 -35.325 ;
        RECT 54.885 -36.475 55.215 -35.325 ;
        RECT 55.450 -35.450 57.100 -35.325 ;
        RECT 58.605 -35.825 58.935 -35.325 ;
        RECT 59.530 -35.785 59.795 -35.325 ;
        RECT 61.700 -36.125 61.870 -35.325 ;
        RECT 63.580 -35.825 63.895 -35.325 ;
        RECT 64.640 -36.335 64.810 -35.325 ;
        RECT 65.480 -36.240 65.655 -35.325 ;
        RECT 66.515 -36.465 66.730 -35.325 ;
        RECT 67.405 -36.465 67.655 -35.325 ;
        RECT 78.700 -35.715 79.030 -34.955 ;
        RECT 68.100 -36.450 68.600 -36.050 ;
        RECT 79.630 -36.105 79.890 -34.955 ;
        RECT 80.600 -35.730 81.000 -35.230 ;
        RECT 82.095 -35.455 82.425 -34.955 ;
        RECT 83.035 -35.455 83.365 -34.955 ;
        RECT 85.010 -35.335 85.390 -34.955 ;
        RECT 85.910 -35.335 86.240 -34.955 ;
        RECT 87.520 -35.335 87.940 -34.955 ;
        RECT 88.610 -35.645 88.940 -34.955 ;
        RECT 90.060 -35.755 90.345 -34.955 ;
        RECT 93.610 -35.715 93.940 -34.955 ;
        RECT 94.540 -35.130 97.350 -34.955 ;
        RECT 94.540 -36.105 94.800 -35.130 ;
        RECT 79.500 -39.995 86.650 -39.980 ;
        RECT 78.290 -40.165 86.650 -39.995 ;
        RECT 77.600 -40.780 78.000 -40.280 ;
        RECT 78.415 -41.305 78.645 -40.165 ;
        RECT 79.315 -40.330 86.650 -40.165 ;
        RECT 79.315 -41.305 79.525 -40.330 ;
        RECT 86.300 -40.465 86.650 -40.330 ;
        RECT 86.300 -40.635 89.520 -40.465 ;
        RECT 90.880 -40.480 92.720 -40.465 ;
        RECT 97.000 -40.480 97.350 -35.130 ;
        RECT 90.880 -40.635 97.350 -40.480 ;
        RECT 87.355 -41.485 87.525 -40.635 ;
        RECT 88.195 -41.145 88.365 -40.635 ;
        RECT 90.050 -41.530 90.450 -41.030 ;
        RECT 91.440 -41.395 91.770 -40.635 ;
        RECT 92.370 -40.830 97.350 -40.635 ;
        RECT 92.370 -41.785 92.630 -40.830 ;
        RECT 20.975 -42.550 21.145 -41.990 ;
        RECT 20.215 -42.880 21.145 -42.550 ;
        RECT 66.800 -42.655 68.150 -42.500 ;
        RECT 54.890 -42.825 57.190 -42.655 ;
        RECT 59.490 -42.825 68.150 -42.655 ;
        RECT 20.975 -43.480 21.145 -42.880 ;
        RECT 19.825 -43.740 21.145 -43.480 ;
        RECT 52.950 -43.550 53.350 -43.050 ;
        RECT 20.975 -43.830 21.145 -43.740 ;
        RECT 55.020 -43.965 55.285 -42.825 ;
        RECT 55.955 -43.625 56.125 -42.825 ;
        RECT 56.795 -43.285 57.005 -42.825 ;
        RECT 60.005 -43.325 60.335 -42.825 ;
        RECT 60.930 -43.285 61.195 -42.825 ;
        RECT 63.100 -43.625 63.270 -42.825 ;
        RECT 64.980 -43.325 65.295 -42.825 ;
        RECT 66.035 -43.835 66.205 -42.825 ;
        RECT 66.800 -42.850 68.150 -42.825 ;
        RECT 20.000 -44.450 20.500 -44.050 ;
        RECT 20.975 -45.415 21.145 -45.290 ;
        RECT 19.835 -45.645 21.145 -45.415 ;
        RECT 20.975 -46.315 21.145 -45.645 ;
        RECT 19.835 -46.525 21.145 -46.315 ;
        RECT 20.975 -46.670 21.145 -46.525 ;
        RECT 67.750 -46.600 68.150 -42.850 ;
        RECT 55.450 -46.855 57.100 -46.700 ;
        RECT 52.690 -47.025 57.100 -46.855 ;
        RECT 58.090 -47.025 67.750 -46.855 ;
        RECT 51.950 -47.800 52.350 -47.300 ;
        RECT 53.285 -47.825 53.525 -47.025 ;
        RECT 54.045 -47.825 54.375 -47.025 ;
        RECT 54.885 -48.175 55.215 -47.025 ;
        RECT 55.450 -47.150 57.100 -47.025 ;
        RECT 58.605 -47.525 58.935 -47.025 ;
        RECT 59.530 -47.485 59.795 -47.025 ;
        RECT 61.700 -47.825 61.870 -47.025 ;
        RECT 63.580 -47.525 63.895 -47.025 ;
        RECT 64.640 -48.035 64.810 -47.025 ;
        RECT 65.480 -47.940 65.655 -47.025 ;
        RECT 66.515 -48.165 66.730 -47.025 ;
        RECT 67.405 -48.165 67.655 -47.025 ;
        RECT 68.100 -48.150 68.600 -47.750 ;
        RECT 79.295 -47.875 79.505 -46.735 ;
        RECT 80.175 -47.875 80.405 -46.735 ;
        RECT 81.000 -47.480 81.400 -46.980 ;
        RECT 82.515 -47.875 82.800 -47.075 ;
        RECT 83.920 -47.875 84.250 -47.185 ;
        RECT 84.920 -47.875 85.340 -47.495 ;
        RECT 86.620 -47.875 86.950 -47.495 ;
        RECT 87.470 -47.875 87.850 -47.495 ;
        RECT 89.495 -47.875 89.825 -47.375 ;
        RECT 90.435 -47.875 90.765 -47.375 ;
        RECT 93.300 -47.875 93.560 -46.725 ;
        RECT 94.160 -47.875 94.490 -47.115 ;
        RECT 97.000 -47.830 97.350 -40.830 ;
        RECT 95.000 -47.875 97.350 -47.830 ;
        RECT 79.150 -48.045 80.530 -47.875 ;
        RECT 81.620 -48.045 91.280 -47.875 ;
        RECT 93.210 -48.045 97.350 -47.875 ;
        RECT 95.000 -48.180 97.350 -48.045 ;
      LAYER met1 ;
        RECT -13.700 20.050 -12.400 21.350 ;
        RECT 15.450 20.250 19.650 20.750 ;
        RECT 15.550 19.550 16.050 20.250 ;
        RECT 15.540 19.070 17.840 19.550 ;
        RECT 18.100 18.450 18.500 20.250 ;
        RECT 17.350 18.050 17.950 18.350 ;
        RECT 19.150 18.050 19.650 20.250 ;
        RECT 17.350 17.750 19.650 18.050 ;
        RECT 74.650 -7.980 104.420 -7.500 ;
        RECT 74.650 -8.000 80.050 -7.980 ;
        RECT 83.600 -8.000 84.100 -7.980 ;
        RECT 87.700 -8.000 88.200 -7.980 ;
        RECT 91.800 -8.000 92.550 -7.980 ;
        RECT 96.200 -8.000 96.650 -7.980 ;
        RECT 100.300 -8.000 100.750 -7.980 ;
        RECT -15.210 -13.060 1.540 -12.580 ;
        RECT -13.400 -13.080 -11.700 -13.060 ;
        RECT -2.150 -13.080 -0.300 -13.060 ;
        RECT -12.750 -13.680 -12.350 -13.080 ;
        RECT 3.650 -13.150 6.200 -12.750 ;
        RECT 28.900 -15.550 31.840 -15.100 ;
        RECT 28.900 -16.270 29.200 -15.550 ;
        RECT 29.540 -15.580 31.840 -15.550 ;
        RECT 32.700 -16.750 33.150 -15.100 ;
        RECT 31.500 -17.100 33.150 -16.750 ;
        RECT -15.750 -17.790 -15.000 -17.780 ;
        RECT -15.750 -18.270 -13.680 -17.790 ;
        RECT -3.850 -18.260 -2.450 -18.230 ;
        RECT -15.750 -18.280 -15.000 -18.270 ;
        RECT -15.750 -18.730 -15.350 -18.280 ;
        RECT -7.050 -18.730 -0.630 -18.260 ;
        RECT -7.050 -18.740 -3.830 -18.730 ;
        RECT -3.300 -19.480 -2.900 -18.730 ;
        RECT -2.470 -18.740 -0.630 -18.730 ;
        RECT -14.200 -25.680 -12.820 -25.670 ;
        RECT -12.350 -25.680 -11.950 -24.930 ;
        RECT -11.730 -25.680 -2.070 -25.670 ;
        RECT -0.140 -25.680 1.700 -25.670 ;
        RECT -14.200 -26.130 1.700 -25.680 ;
        RECT -14.200 -26.150 -12.820 -26.130 ;
        RECT -11.730 -26.150 -2.070 -26.130 ;
        RECT -0.140 -26.150 1.700 -26.130 ;
        RECT 49.000 -28.100 49.550 -27.300 ;
        RECT 52.850 -27.375 55.400 -27.300 ;
        RECT 74.650 -27.375 75.150 -8.000 ;
        RECT 77.250 -11.500 77.750 -8.000 ;
        RECT 92.050 -8.650 92.450 -8.000 ;
        RECT 77.250 -11.980 81.780 -11.500 ;
        RECT 83.740 -11.980 97.020 -11.500 ;
        RECT 77.250 -12.000 80.050 -11.980 ;
        RECT 91.100 -12.000 93.000 -11.980 ;
        RECT 94.350 -12.000 95.650 -11.980 ;
        RECT 82.200 -12.650 82.600 -12.150 ;
        RECT 52.850 -27.800 78.600 -27.375 ;
        RECT 54.975 -27.825 78.600 -27.800 ;
        RECT 47.140 -28.550 49.550 -28.100 ;
        RECT 47.140 -28.580 48.980 -28.550 ;
        RECT 49.250 -29.500 49.550 -28.550 ;
        RECT 54.890 -31.280 66.850 -30.800 ;
        RECT 57.150 -31.300 59.600 -31.280 ;
        RECT 51.100 -31.850 53.350 -31.350 ;
        RECT 51.100 -35.600 51.600 -31.850 ;
        RECT 67.750 -35.000 68.150 -34.500 ;
        RECT 78.150 -34.630 78.600 -27.825 ;
        RECT 52.690 -35.480 55.450 -35.000 ;
        RECT 56.600 -35.450 68.150 -35.000 ;
        RECT 78.140 -35.110 94.890 -34.630 ;
        RECT 79.950 -35.130 81.650 -35.110 ;
        RECT 91.200 -35.130 93.050 -35.110 ;
        RECT 58.090 -35.480 68.150 -35.450 ;
        RECT 67.750 -35.500 68.150 -35.480 ;
        RECT 51.100 -36.100 52.350 -35.600 ;
        RECT 80.600 -35.730 81.000 -35.130 ;
        RECT 68.100 -36.450 68.600 -36.050 ;
        RECT 77.600 -39.840 78.350 -39.830 ;
        RECT 77.600 -40.320 79.670 -39.840 ;
        RECT 89.500 -40.310 90.900 -40.280 ;
        RECT 77.600 -40.330 78.350 -40.320 ;
        RECT 77.600 -40.780 78.000 -40.330 ;
        RECT 86.300 -40.780 92.720 -40.310 ;
        RECT 86.300 -40.790 89.520 -40.780 ;
        RECT 20.800 -42.000 21.300 -40.950 ;
        RECT 90.050 -41.530 90.450 -40.780 ;
        RECT 90.880 -40.790 92.720 -40.780 ;
        RECT 20.820 -43.800 21.300 -42.000 ;
        RECT 54.890 -42.980 66.850 -42.500 ;
        RECT 57.150 -43.000 59.600 -42.980 ;
        RECT 45.750 -43.550 53.350 -43.050 ;
        RECT 20.800 -44.050 21.300 -43.800 ;
        RECT 20.000 -44.450 21.300 -44.050 ;
        RECT 20.800 -45.300 21.300 -44.450 ;
        RECT 20.820 -46.670 21.300 -45.300 ;
        RECT 51.100 -46.700 51.600 -43.550 ;
        RECT 67.750 -46.700 68.150 -46.200 ;
        RECT 51.100 -47.150 55.450 -46.700 ;
        RECT 56.600 -47.150 68.150 -46.700 ;
        RECT 51.100 -47.300 51.600 -47.150 ;
        RECT 52.690 -47.180 55.450 -47.150 ;
        RECT 58.090 -47.180 68.150 -47.150 ;
        RECT 67.750 -47.200 68.150 -47.180 ;
        RECT 51.100 -47.800 52.350 -47.300 ;
        RECT 79.150 -47.730 80.530 -47.720 ;
        RECT 81.000 -47.730 81.400 -46.980 ;
        RECT 81.620 -47.730 91.280 -47.720 ;
        RECT 93.210 -47.730 95.050 -47.720 ;
        RECT 68.100 -48.150 68.600 -47.750 ;
        RECT 79.150 -48.180 95.050 -47.730 ;
        RECT 79.150 -48.200 80.530 -48.180 ;
        RECT 81.620 -48.200 91.280 -48.180 ;
        RECT 93.210 -48.200 95.050 -48.180 ;
      LAYER met2 ;
        RECT -13.700 20.050 -12.400 21.350 ;
        RECT -13.525 -0.825 -12.575 20.050 ;
        RECT -13.525 -1.775 10.450 -0.825 ;
        RECT 9.500 -12.750 10.450 -1.775 ;
        RECT 3.650 -13.150 10.450 -12.750 ;
        RECT 9.500 -15.100 10.450 -13.150 ;
        RECT 9.500 -15.550 33.150 -15.100 ;
        RECT 9.500 -27.300 10.450 -15.550 ;
        RECT 9.500 -27.750 55.400 -27.300 ;
        RECT 9.500 -33.525 10.450 -27.750 ;
        RECT 20.800 -41.450 21.300 -27.750 ;
        RECT 45.750 -43.550 46.250 -27.750 ;
        RECT 52.850 -27.800 55.400 -27.750 ;
    END
  END VCCD
  PIN ENB
    ANTENNAGATEAREA 1.437000 ;
    PORT
      LAYER li1 ;
        RECT 15.625 18.250 16.085 18.315 ;
        RECT -22.350 17.950 16.085 18.250 ;
        RECT -22.350 -8.750 -22.050 17.950 ;
        RECT 15.625 17.585 16.085 17.950 ;
        RECT -22.350 -9.150 7.150 -8.750 ;
        RECT -22.350 -58.400 -22.050 -9.150 ;
        RECT 6.750 -16.750 7.150 -9.150 ;
        RECT 6.750 -17.150 27.850 -16.750 ;
        RECT 29.625 -17.065 30.085 -16.335 ;
        RECT -14.955 -19.675 -14.625 -19.425 ;
        RECT 76.400 -58.400 76.900 -41.350 ;
        RECT 78.395 -41.725 78.725 -41.475 ;
        RECT -22.350 -58.900 76.900 -58.400 ;
      LAYER met1 ;
        RECT 27.500 -16.800 27.850 -16.750 ;
        RECT 29.600 -16.800 30.100 -16.550 ;
        RECT 27.500 -17.100 30.100 -16.800 ;
        RECT 27.500 -17.150 27.850 -17.100 ;
        RECT -22.350 -19.380 -15.800 -19.350 ;
        RECT -22.350 -19.730 -14.600 -19.380 ;
        RECT -22.350 -19.750 -15.800 -19.730 ;
        RECT 76.400 -41.430 76.900 -41.350 ;
        RECT 76.400 -41.780 78.750 -41.430 ;
        RECT 76.400 -41.850 76.900 -41.780 ;
    END
  END ENB
  PIN GND
    ANTENNADIFFAREA 61.479050 ;
    PORT
      LAYER pwell ;
        RECT -7.100 26.800 82.900 31.600 ;
        RECT 16.030 17.600 17.835 17.605 ;
        RECT 16.030 17.375 18.750 17.600 ;
        RECT 15.545 16.700 18.750 17.375 ;
        RECT 15.545 16.695 17.835 16.700 ;
        RECT 15.690 16.505 15.860 16.695 ;
        RECT 22.900 11.850 82.900 16.650 ;
        RECT 21.500 -12.450 64.700 -9.650 ;
        RECT 79.750 -10.400 104.650 -9.400 ;
        RECT 80.085 -10.545 80.255 -10.400 ;
        RECT 84.185 -10.545 84.355 -10.400 ;
        RECT 88.285 -10.545 88.455 -10.400 ;
        RECT 92.685 -10.545 92.855 -10.400 ;
        RECT 96.785 -10.545 96.955 -10.400 ;
        RECT 100.885 -10.545 101.055 -10.400 ;
        RECT 79.750 -14.400 97.250 -13.400 ;
        RECT -14.720 -14.730 -13.375 -14.525 ;
        RECT -16.000 -14.755 -15.150 -14.730 ;
        RECT -14.720 -14.755 -11.750 -14.730 ;
        RECT -10.405 -14.755 -9.485 -14.535 ;
        RECT -3.405 -14.635 -2.485 -14.525 ;
        RECT -4.820 -14.730 -2.485 -14.635 ;
        RECT -4.820 -14.755 -0.250 -14.730 ;
        RECT 0.190 -14.755 1.535 -14.525 ;
        RECT 80.085 -14.545 80.255 -14.400 ;
        RECT 83.885 -14.545 84.055 -14.400 ;
        RECT 93.130 -14.545 93.300 -14.400 ;
        RECT 95.785 -14.545 95.955 -14.400 ;
        RECT -16.000 -15.430 1.535 -14.755 ;
        RECT -15.205 -15.435 -13.375 -15.430 ;
        RECT -11.765 -15.435 -2.485 -15.430 ;
        RECT -0.295 -15.435 1.535 -15.430 ;
        RECT -15.065 -15.625 -14.895 -15.435 ;
        RECT -11.625 -15.625 -11.455 -15.435 ;
        RECT -0.155 -15.625 0.015 -15.435 ;
        RECT 30.030 -17.275 31.835 -17.045 ;
        RECT 29.545 -17.280 31.835 -17.275 ;
        RECT 28.880 -17.955 31.835 -17.280 ;
        RECT 28.880 -17.960 29.550 -17.955 ;
        RECT 29.690 -18.145 29.860 -17.955 ;
        RECT -15.950 -19.735 -15.000 -19.730 ;
        RECT -15.950 -20.630 -13.695 -19.735 ;
        RECT -15.045 -20.645 -13.695 -20.630 ;
        RECT -7.005 -20.430 -3.835 -20.205 ;
        RECT -7.005 -20.435 -2.450 -20.430 ;
        RECT -1.980 -20.435 -0.635 -20.205 ;
        RECT -14.915 -20.835 -14.745 -20.645 ;
        RECT -7.005 -21.115 -0.635 -20.435 ;
        RECT 35.950 -20.650 64.750 -17.850 ;
        RECT -6.905 -21.305 -6.735 -21.115 ;
        RECT -3.850 -21.130 -2.450 -21.115 ;
        RECT -2.325 -21.305 -2.155 -21.115 ;
        RECT -13.135 -23.295 -12.965 -23.105 ;
        RECT -12.850 -23.295 -11.350 -23.280 ;
        RECT -2.385 -23.295 -2.215 -23.105 ;
        RECT -2.100 -23.295 -0.100 -23.280 ;
        RECT 1.385 -23.295 1.555 -23.105 ;
        RECT -14.185 -23.975 1.695 -23.295 ;
        RECT -14.185 -24.095 -9.020 -23.975 ;
        RECT -14.185 -24.205 -10.435 -24.095 ;
        RECT -4.355 -24.195 -3.435 -23.975 ;
        RECT -2.100 -23.980 1.210 -23.975 ;
        RECT -0.135 -24.205 1.210 -23.980 ;
        RECT -12.850 -24.230 -11.350 -24.205 ;
        RECT 47.630 -30.050 48.975 -30.045 ;
        RECT 47.630 -30.275 49.800 -30.050 ;
        RECT 47.145 -30.950 49.800 -30.275 ;
        RECT 47.145 -30.955 48.975 -30.950 ;
        RECT 47.285 -31.145 47.455 -30.955 ;
        RECT 52.650 -32.745 55.000 -32.700 ;
        RECT 52.650 -32.950 57.135 -32.745 ;
        RECT 52.650 -32.975 59.550 -32.950 ;
        RECT 63.010 -32.975 63.920 -32.755 ;
        RECT 65.455 -32.975 66.805 -32.745 ;
        RECT 52.650 -33.655 66.805 -32.975 ;
        RECT 52.650 -33.700 55.000 -33.655 ;
        RECT 55.035 -33.845 55.205 -33.655 ;
        RECT 57.100 -33.700 59.550 -33.655 ;
        RECT 59.635 -33.845 59.805 -33.655 ;
        RECT 78.630 -36.780 79.975 -36.575 ;
        RECT 77.350 -36.805 78.200 -36.780 ;
        RECT 78.630 -36.805 81.600 -36.780 ;
        RECT 82.945 -36.805 83.865 -36.585 ;
        RECT 89.945 -36.685 90.865 -36.575 ;
        RECT 88.530 -36.780 90.865 -36.685 ;
        RECT 88.530 -36.805 93.100 -36.780 ;
        RECT 93.540 -36.805 94.885 -36.575 ;
        RECT 52.695 -36.950 55.305 -36.945 ;
        RECT 51.650 -37.150 55.305 -36.950 ;
        RECT 51.650 -37.175 58.150 -37.150 ;
        RECT 61.610 -37.175 62.520 -36.955 ;
        RECT 64.060 -37.175 67.745 -36.945 ;
        RECT 51.650 -37.855 67.745 -37.175 ;
        RECT 77.350 -37.480 94.885 -36.805 ;
        RECT 78.145 -37.485 79.975 -37.480 ;
        RECT 81.585 -37.485 90.865 -37.480 ;
        RECT 93.055 -37.485 94.885 -37.480 ;
        RECT 78.285 -37.675 78.455 -37.485 ;
        RECT 81.725 -37.675 81.895 -37.485 ;
        RECT 93.195 -37.675 93.365 -37.485 ;
        RECT 51.650 -38.200 52.750 -37.855 ;
        RECT 52.840 -38.045 53.010 -37.855 ;
        RECT 55.300 -37.900 58.150 -37.855 ;
        RECT 58.235 -38.045 58.405 -37.855 ;
        RECT 18.445 -42.135 19.125 -41.995 ;
        RECT 18.255 -42.305 19.125 -42.135 ;
        RECT 18.445 -42.480 19.125 -42.305 ;
        RECT 29.650 -42.350 32.950 -39.550 ;
        RECT 34.200 -42.350 37.500 -39.550 ;
        RECT 77.400 -41.785 78.350 -41.780 ;
        RECT 18.445 -43.825 19.355 -42.480 ;
        RECT 77.400 -42.680 79.655 -41.785 ;
        RECT 78.305 -42.695 79.655 -42.680 ;
        RECT 86.345 -42.480 89.515 -42.255 ;
        RECT 86.345 -42.485 90.900 -42.480 ;
        RECT 91.370 -42.485 92.715 -42.255 ;
        RECT 78.435 -42.885 78.605 -42.695 ;
        RECT 86.345 -43.165 92.715 -42.485 ;
        RECT 86.445 -43.355 86.615 -43.165 ;
        RECT 89.500 -43.180 90.900 -43.165 ;
        RECT 91.025 -43.355 91.195 -43.165 ;
        RECT 18.450 -45.305 19.350 -43.825 ;
        RECT 52.650 -44.445 55.000 -44.400 ;
        RECT 52.650 -44.650 57.135 -44.445 ;
        RECT 52.650 -44.675 59.550 -44.650 ;
        RECT 63.010 -44.675 63.920 -44.455 ;
        RECT 65.455 -44.675 66.805 -44.445 ;
        RECT 18.445 -45.435 19.355 -45.305 ;
        RECT 52.650 -45.355 66.805 -44.675 ;
        RECT 80.215 -45.345 80.385 -45.155 ;
        RECT 80.500 -45.345 82.000 -45.330 ;
        RECT 90.965 -45.345 91.135 -45.155 ;
        RECT 91.250 -45.345 93.250 -45.330 ;
        RECT 94.735 -45.345 94.905 -45.155 ;
        RECT 52.650 -45.400 55.000 -45.355 ;
        RECT 18.255 -45.605 19.355 -45.435 ;
        RECT 55.035 -45.545 55.205 -45.355 ;
        RECT 57.100 -45.400 59.550 -45.355 ;
        RECT 59.635 -45.545 59.805 -45.355 ;
        RECT 18.445 -46.655 19.355 -45.605 ;
        RECT 79.165 -46.025 95.045 -45.345 ;
        RECT 79.165 -46.145 84.330 -46.025 ;
        RECT 79.165 -46.255 82.915 -46.145 ;
        RECT 88.995 -46.245 89.915 -46.025 ;
        RECT 91.250 -46.030 94.560 -46.025 ;
        RECT 93.215 -46.255 94.560 -46.030 ;
        RECT 80.500 -46.280 82.000 -46.255 ;
        RECT 27.100 -50.350 41.480 -48.340 ;
        RECT 52.695 -48.650 55.305 -48.645 ;
        RECT 51.650 -48.850 55.305 -48.650 ;
        RECT 51.650 -48.875 58.150 -48.850 ;
        RECT 61.610 -48.875 62.520 -48.655 ;
        RECT 64.060 -48.875 67.745 -48.645 ;
        RECT 51.650 -49.555 67.745 -48.875 ;
        RECT 51.650 -49.900 52.750 -49.555 ;
        RECT 52.840 -49.745 53.010 -49.555 ;
        RECT 55.300 -49.600 58.150 -49.555 ;
        RECT 58.235 -49.745 58.405 -49.555 ;
      LAYER li1 ;
        RECT -6.900 27.150 -6.500 27.650 ;
        RECT 2.600 27.150 3.000 27.650 ;
        RECT 8.050 27.150 8.450 27.650 ;
        RECT 13.500 27.150 13.900 27.650 ;
        RECT 23.100 27.150 23.500 27.650 ;
        RECT 32.600 27.150 33.000 27.650 ;
        RECT 38.050 27.150 38.450 27.650 ;
        RECT 43.500 27.150 43.900 27.650 ;
        RECT 53.100 27.150 53.500 27.650 ;
        RECT 62.600 27.150 63.000 27.650 ;
        RECT 68.050 27.150 68.450 27.650 ;
        RECT 73.500 27.150 73.900 27.650 ;
        RECT 31.000 21.250 31.170 21.330 ;
        RECT 29.185 20.930 31.170 21.250 ;
        RECT 31.000 20.850 31.170 20.930 ;
        RECT 16.055 16.675 16.990 17.075 ;
        RECT 18.100 16.950 18.500 17.450 ;
        RECT 15.540 16.505 17.840 16.675 ;
        RECT 31.900 15.800 32.300 16.300 ;
        RECT 37.350 15.800 37.750 16.300 ;
        RECT 42.800 15.800 43.200 16.300 ;
        RECT 52.300 15.800 52.700 16.300 ;
        RECT 61.900 15.800 62.300 16.300 ;
        RECT 67.350 15.800 67.750 16.300 ;
        RECT 72.800 15.800 73.200 16.300 ;
        RECT 82.300 15.800 82.700 16.300 ;
        RECT 21.700 -12.100 22.100 -11.600 ;
        RECT 22.400 -12.950 22.800 -10.050 ;
        RECT 25.200 -12.950 25.600 -10.050 ;
        RECT 26.000 -12.100 26.400 -11.600 ;
        RECT 26.700 -12.950 27.100 -10.050 ;
        RECT 28.900 -12.100 29.300 -11.600 ;
        RECT 29.600 -12.950 30.000 -10.050 ;
        RECT 31.800 -12.100 32.200 -11.600 ;
        RECT 32.500 -12.950 32.900 -10.050 ;
        RECT 35.300 -12.950 35.700 -10.050 ;
        RECT 36.100 -12.100 36.500 -11.600 ;
        RECT 36.800 -12.950 37.200 -10.050 ;
        RECT 39.600 -12.950 40.000 -10.050 ;
        RECT 40.400 -12.100 40.800 -11.600 ;
        RECT 41.100 -12.950 41.500 -10.050 ;
        RECT 43.300 -12.100 43.700 -11.600 ;
        RECT 44.000 -12.950 44.400 -10.050 ;
        RECT 46.200 -12.100 46.600 -11.600 ;
        RECT 46.900 -12.950 47.300 -10.050 ;
        RECT 49.700 -12.950 50.100 -10.050 ;
        RECT 50.500 -12.100 50.900 -11.600 ;
        RECT 51.200 -12.950 51.600 -10.050 ;
        RECT 54.000 -12.950 54.400 -10.050 ;
        RECT 54.800 -12.100 55.200 -11.600 ;
        RECT 55.500 -12.950 55.900 -10.050 ;
        RECT 57.700 -12.100 58.100 -11.600 ;
        RECT 58.400 -12.950 58.800 -10.050 ;
        RECT 60.600 -12.100 61.000 -11.600 ;
        RECT 61.300 -12.950 61.700 -10.050 ;
        RECT 64.100 -12.950 64.500 -10.050 ;
        RECT 80.595 -10.375 80.865 -9.915 ;
        RECT 82.655 -10.375 82.980 -9.915 ;
        RECT 84.695 -10.375 84.965 -9.915 ;
        RECT 86.755 -10.375 87.080 -9.915 ;
        RECT 88.795 -10.375 89.065 -9.915 ;
        RECT 90.855 -10.375 91.180 -9.915 ;
        RECT 92.000 -10.210 92.310 -9.710 ;
        RECT 93.195 -10.375 93.465 -9.915 ;
        RECT 95.255 -10.375 95.580 -9.915 ;
        RECT 97.295 -10.375 97.565 -9.915 ;
        RECT 99.355 -10.375 99.680 -9.915 ;
        RECT 101.395 -10.375 101.665 -9.915 ;
        RECT 103.455 -10.375 103.780 -9.915 ;
        RECT 79.940 -10.545 83.620 -10.375 ;
        RECT 84.040 -10.545 87.720 -10.375 ;
        RECT 88.140 -10.545 91.820 -10.375 ;
        RECT 92.540 -10.545 96.220 -10.375 ;
        RECT 96.640 -10.545 100.320 -10.375 ;
        RECT 100.740 -10.545 104.420 -10.375 ;
        RECT 22.400 -13.350 64.500 -12.950 ;
        RECT -15.800 -15.280 -15.400 -14.780 ;
        RECT -14.650 -15.455 -14.320 -15.075 ;
        RECT -13.720 -15.280 -13.460 -14.615 ;
        RECT -13.720 -15.455 -11.750 -15.280 ;
        RECT -11.255 -15.455 -10.925 -15.075 ;
        RECT -10.315 -15.455 -9.985 -15.075 ;
        RECT -8.160 -15.455 -7.750 -15.015 ;
        RECT -7.010 -15.455 -6.690 -14.995 ;
        RECT -5.080 -15.455 -4.420 -14.975 ;
        RECT -3.290 -15.455 -3.005 -14.995 ;
        RECT -2.150 -15.455 -0.300 -15.330 ;
        RECT 0.260 -15.455 0.590 -15.075 ;
        RECT 1.190 -15.455 1.450 -14.615 ;
        RECT -15.210 -15.625 1.540 -15.455 ;
        RECT -13.500 -15.780 -11.750 -15.625 ;
        RECT -2.150 -15.780 -0.300 -15.625 ;
        RECT 36.150 -16.950 36.550 -13.350 ;
        RECT 63.450 -16.950 63.850 -13.350 ;
        RECT 80.500 -14.375 80.830 -13.995 ;
        RECT 81.430 -14.375 81.690 -13.535 ;
        RECT 81.950 -14.100 82.350 -13.600 ;
        RECT 84.255 -14.375 84.585 -13.995 ;
        RECT 85.195 -14.375 85.445 -13.915 ;
        RECT 87.140 -14.375 87.510 -13.875 ;
        RECT 89.325 -14.375 89.535 -13.845 ;
        RECT 90.295 -14.375 90.465 -13.765 ;
        RECT 93.075 -14.375 93.385 -13.575 ;
        RECT 95.765 -14.375 95.995 -13.555 ;
        RECT 96.665 -14.375 96.875 -13.555 ;
        RECT 79.940 -14.545 81.780 -14.375 ;
        RECT 83.740 -14.545 91.100 -14.375 ;
        RECT 92.990 -14.545 94.370 -14.375 ;
        RECT 95.640 -14.545 97.020 -14.375 ;
        RECT 35.100 -17.350 63.850 -16.950 ;
        RECT 28.950 -18.400 29.300 -17.350 ;
        RECT 30.055 -17.975 30.990 -17.575 ;
        RECT 29.540 -18.145 31.840 -17.975 ;
        RECT 29.550 -18.400 29.900 -18.145 ;
        RECT 28.950 -18.750 29.900 -18.400 ;
        RECT -15.750 -20.480 -15.350 -19.980 ;
        RECT -14.935 -20.665 -14.705 -19.845 ;
        RECT -14.035 -20.480 -13.825 -19.845 ;
        RECT -14.035 -20.665 -9.150 -20.480 ;
        RECT -15.060 -20.830 -9.150 -20.665 ;
        RECT -15.060 -20.835 -13.680 -20.830 ;
        RECT -9.500 -21.030 -9.150 -20.830 ;
        RECT -6.915 -21.030 -6.585 -20.745 ;
        RECT -9.500 -21.135 -6.585 -21.030 ;
        RECT -6.075 -21.135 -5.745 -20.745 ;
        RECT -4.205 -21.135 -3.915 -20.300 ;
        RECT -3.400 -20.980 -2.900 -20.580 ;
        RECT -1.910 -21.135 -1.580 -20.755 ;
        RECT -0.980 -21.135 -0.720 -20.295 ;
        RECT 28.950 -20.600 29.450 -18.750 ;
        RECT 35.100 -20.600 35.500 -17.350 ;
        RECT 36.150 -20.250 36.550 -17.350 ;
        RECT 38.950 -20.250 39.350 -17.350 ;
        RECT 39.650 -18.700 40.050 -18.200 ;
        RECT 41.850 -20.250 42.250 -17.350 ;
        RECT 42.550 -18.700 42.950 -18.200 ;
        RECT 44.750 -20.250 45.150 -17.350 ;
        RECT 45.450 -18.700 45.850 -18.200 ;
        RECT 46.250 -20.250 46.650 -17.350 ;
        RECT 49.050 -20.250 49.450 -17.350 ;
        RECT 49.750 -18.700 50.150 -18.200 ;
        RECT 50.550 -20.250 50.950 -17.350 ;
        RECT 53.350 -20.250 53.750 -17.350 ;
        RECT 54.050 -18.700 54.450 -18.200 ;
        RECT 56.250 -20.250 56.650 -17.350 ;
        RECT 56.950 -18.700 57.350 -18.200 ;
        RECT 59.150 -20.250 59.550 -17.350 ;
        RECT 59.850 -18.700 60.250 -18.200 ;
        RECT 60.650 -20.250 61.050 -17.350 ;
        RECT 63.450 -20.250 63.850 -17.350 ;
        RECT 64.150 -18.700 64.550 -18.200 ;
        RECT 28.950 -21.000 35.500 -20.600 ;
        RECT -9.500 -21.305 -3.830 -21.135 ;
        RECT -2.470 -21.305 -0.630 -21.135 ;
        RECT -9.500 -21.380 -6.850 -21.305 ;
        RECT -12.950 -23.105 -11.650 -22.980 ;
        RECT -9.500 -23.105 -9.150 -21.380 ;
        RECT -2.100 -23.105 0.050 -23.080 ;
        RECT -14.200 -23.275 1.700 -23.105 ;
        RECT -14.055 -24.095 -13.845 -23.275 ;
        RECT -13.175 -23.430 -11.650 -23.275 ;
        RECT -13.175 -24.095 -12.945 -23.430 ;
        RECT -10.835 -23.735 -10.550 -23.275 ;
        RECT -9.420 -23.755 -8.760 -23.275 ;
        RECT -7.150 -23.735 -6.830 -23.275 ;
        RECT -6.090 -23.715 -5.680 -23.275 ;
        RECT -3.855 -23.655 -3.525 -23.275 ;
        RECT -2.915 -23.655 -2.585 -23.275 ;
        RECT -2.100 -23.430 0.210 -23.275 ;
        RECT -1.000 -23.830 -0.500 -23.430 ;
        RECT -0.050 -24.115 0.210 -23.430 ;
        RECT 0.810 -23.655 1.140 -23.275 ;
        RECT 28.950 -29.550 29.450 -21.000 ;
        RECT 47.700 -30.975 48.030 -30.595 ;
        RECT 48.630 -30.975 48.890 -30.135 ;
        RECT 47.140 -31.145 48.980 -30.975 ;
        RECT 48.550 -31.800 48.950 -31.145 ;
        RECT 49.250 -31.800 49.550 -30.250 ;
        RECT 48.550 -32.100 49.550 -31.800 ;
        RECT 48.550 -33.000 48.950 -32.100 ;
        RECT 48.550 -33.500 53.350 -33.000 ;
        RECT 48.550 -33.700 49.050 -33.500 ;
        RECT 55.020 -33.650 55.285 -33.215 ;
        RECT 55.020 -33.675 55.300 -33.650 ;
        RECT 55.955 -33.675 56.125 -33.215 ;
        RECT 56.795 -33.675 57.045 -33.210 ;
        RECT 60.005 -33.675 60.335 -33.295 ;
        RECT 60.945 -33.675 61.195 -33.215 ;
        RECT 62.890 -33.675 63.260 -33.175 ;
        RECT 65.075 -33.675 65.285 -33.145 ;
        RECT 66.045 -33.675 66.215 -33.065 ;
        RECT 54.890 -33.700 57.190 -33.675 ;
        RECT 48.550 -33.845 57.190 -33.700 ;
        RECT 59.490 -33.845 66.850 -33.675 ;
        RECT 48.550 -34.100 55.300 -33.845 ;
        RECT 29.850 -40.400 30.250 -39.900 ;
        RECT 18.255 -42.550 18.425 -41.990 ;
        RECT 36.900 -42.000 37.300 -41.500 ;
        RECT 18.255 -42.880 18.805 -42.550 ;
        RECT 18.255 -43.480 18.425 -42.880 ;
        RECT 18.255 -43.740 19.265 -43.480 ;
        RECT 18.255 -43.830 18.425 -43.740 ;
        RECT 18.600 -44.550 19.100 -44.150 ;
        RECT 48.550 -44.700 49.050 -34.100 ;
        RECT 51.950 -37.900 52.350 -37.400 ;
        RECT 53.215 -37.875 53.455 -37.395 ;
        RECT 54.045 -37.875 54.375 -37.395 ;
        RECT 54.885 -37.875 55.215 -37.075 ;
        RECT 55.450 -37.875 58.100 -37.700 ;
        RECT 58.605 -37.875 58.935 -37.495 ;
        RECT 59.545 -37.875 59.795 -37.415 ;
        RECT 61.490 -37.875 61.860 -37.375 ;
        RECT 63.675 -37.875 63.885 -37.345 ;
        RECT 64.650 -37.875 64.820 -37.265 ;
        RECT 65.490 -37.875 65.660 -37.360 ;
        RECT 66.480 -37.875 66.810 -37.135 ;
        RECT 67.405 -37.875 67.655 -37.055 ;
        RECT 77.550 -37.330 77.950 -36.830 ;
        RECT 78.700 -37.505 79.030 -37.125 ;
        RECT 79.630 -37.330 79.890 -36.665 ;
        RECT 79.630 -37.505 81.600 -37.330 ;
        RECT 82.095 -37.505 82.425 -37.125 ;
        RECT 83.035 -37.505 83.365 -37.125 ;
        RECT 85.190 -37.505 85.600 -37.065 ;
        RECT 86.340 -37.505 86.660 -37.045 ;
        RECT 88.270 -37.505 88.930 -37.025 ;
        RECT 90.060 -37.505 90.345 -37.045 ;
        RECT 91.200 -37.505 93.050 -37.380 ;
        RECT 93.610 -37.505 93.940 -37.125 ;
        RECT 94.540 -37.505 94.800 -36.665 ;
        RECT 78.140 -37.675 94.890 -37.505 ;
        RECT 79.850 -37.830 81.600 -37.675 ;
        RECT 91.200 -37.830 93.050 -37.675 ;
        RECT 52.690 -38.045 67.750 -37.875 ;
        RECT 55.450 -38.200 58.100 -38.045 ;
        RECT 77.600 -42.530 78.000 -42.030 ;
        RECT 78.415 -42.715 78.645 -41.895 ;
        RECT 79.315 -42.530 79.525 -41.895 ;
        RECT 79.315 -42.715 84.200 -42.530 ;
        RECT 78.290 -42.880 84.200 -42.715 ;
        RECT 78.290 -42.885 79.670 -42.880 ;
        RECT 83.850 -43.080 84.200 -42.880 ;
        RECT 86.435 -43.080 86.765 -42.795 ;
        RECT 83.850 -43.185 86.765 -43.080 ;
        RECT 87.275 -43.185 87.605 -42.795 ;
        RECT 89.145 -43.185 89.435 -42.350 ;
        RECT 89.950 -43.030 90.450 -42.630 ;
        RECT 91.440 -43.185 91.770 -42.805 ;
        RECT 92.370 -43.185 92.630 -42.345 ;
        RECT 83.850 -43.355 89.520 -43.185 ;
        RECT 90.880 -43.355 92.720 -43.185 ;
        RECT 83.850 -43.430 86.500 -43.355 ;
        RECT 48.550 -45.200 53.350 -44.700 ;
        RECT 18.255 -45.415 18.425 -45.290 ;
        RECT 48.550 -45.400 49.050 -45.200 ;
        RECT 55.020 -45.350 55.285 -44.915 ;
        RECT 55.020 -45.375 55.350 -45.350 ;
        RECT 55.955 -45.375 56.125 -44.915 ;
        RECT 56.795 -45.375 57.045 -44.910 ;
        RECT 60.005 -45.375 60.335 -44.995 ;
        RECT 60.945 -45.375 61.195 -44.915 ;
        RECT 62.890 -45.375 63.260 -44.875 ;
        RECT 65.075 -45.375 65.285 -44.845 ;
        RECT 66.045 -45.375 66.215 -44.765 ;
        RECT 80.400 -45.155 81.700 -45.030 ;
        RECT 83.850 -45.155 84.200 -43.430 ;
        RECT 91.250 -45.155 93.400 -45.130 ;
        RECT 79.150 -45.325 95.050 -45.155 ;
        RECT 54.890 -45.400 57.190 -45.375 ;
        RECT 18.255 -45.645 19.245 -45.415 ;
        RECT 48.550 -45.545 57.190 -45.400 ;
        RECT 59.490 -45.545 66.850 -45.375 ;
        RECT 18.255 -46.315 18.425 -45.645 ;
        RECT 48.550 -45.750 55.350 -45.545 ;
        RECT 18.255 -46.525 19.245 -46.315 ;
        RECT 18.255 -46.670 18.425 -46.525 ;
        RECT 25.400 -47.850 30.250 -47.450 ;
        RECT 27.280 -48.690 41.300 -48.520 ;
        RECT 27.280 -49.850 27.450 -48.690 ;
        RECT 40.550 -49.170 40.850 -49.150 ;
        RECT 38.490 -49.520 40.850 -49.170 ;
        RECT 26.850 -50.000 27.850 -49.850 ;
        RECT 40.550 -50.000 40.850 -49.520 ;
        RECT 41.130 -50.000 41.300 -48.690 ;
        RECT 26.850 -50.170 41.300 -50.000 ;
        RECT 26.850 -54.650 27.850 -50.170 ;
        RECT 48.550 -54.650 49.050 -45.750 ;
        RECT 79.295 -46.145 79.505 -45.325 ;
        RECT 80.175 -45.480 81.700 -45.325 ;
        RECT 80.175 -46.145 80.405 -45.480 ;
        RECT 82.515 -45.785 82.800 -45.325 ;
        RECT 83.930 -45.805 84.590 -45.325 ;
        RECT 86.200 -45.785 86.520 -45.325 ;
        RECT 87.260 -45.765 87.670 -45.325 ;
        RECT 89.495 -45.705 89.825 -45.325 ;
        RECT 90.435 -45.705 90.765 -45.325 ;
        RECT 91.250 -45.480 93.560 -45.325 ;
        RECT 92.350 -45.880 92.850 -45.480 ;
        RECT 93.300 -46.165 93.560 -45.480 ;
        RECT 94.160 -45.705 94.490 -45.325 ;
        RECT 51.950 -49.600 52.350 -49.100 ;
        RECT 53.215 -49.575 53.455 -49.095 ;
        RECT 54.045 -49.575 54.375 -49.095 ;
        RECT 54.885 -49.575 55.215 -48.775 ;
        RECT 55.450 -49.575 58.100 -49.400 ;
        RECT 58.605 -49.575 58.935 -49.195 ;
        RECT 59.545 -49.575 59.795 -49.115 ;
        RECT 61.490 -49.575 61.860 -49.075 ;
        RECT 63.675 -49.575 63.885 -49.045 ;
        RECT 64.650 -49.575 64.820 -48.965 ;
        RECT 65.490 -49.575 65.660 -49.060 ;
        RECT 66.480 -49.575 66.810 -48.835 ;
        RECT 67.405 -49.575 67.655 -48.755 ;
        RECT 52.690 -49.745 67.750 -49.575 ;
        RECT 55.450 -49.900 58.100 -49.745 ;
        RECT 26.850 -55.650 50.200 -54.650 ;
      LAYER met1 ;
        RECT -6.900 24.900 -6.500 27.650 ;
        RECT 2.600 24.900 3.000 27.650 ;
        RECT 8.050 24.900 8.450 27.650 ;
        RECT 13.500 24.900 13.900 27.650 ;
        RECT 23.100 24.900 23.500 27.650 ;
        RECT 32.600 24.900 33.000 27.650 ;
        RECT 38.050 24.900 38.450 27.650 ;
        RECT 43.500 24.900 43.900 27.650 ;
        RECT 53.100 24.900 53.500 27.650 ;
        RECT 62.600 24.900 63.000 27.650 ;
        RECT 68.050 24.900 68.450 27.650 ;
        RECT 73.500 24.900 73.900 27.650 ;
        RECT -6.900 24.400 73.900 24.900 ;
        RECT 18.100 17.300 18.500 17.450 ;
        RECT 21.050 17.300 21.550 24.400 ;
        RECT 31.900 21.350 32.400 24.400 ;
        RECT 31.050 21.280 32.400 21.350 ;
        RECT 29.125 20.900 32.400 21.280 ;
        RECT 31.050 20.800 32.400 20.900 ;
        RECT 18.100 17.000 21.550 17.300 ;
        RECT 18.100 16.950 18.500 17.000 ;
        RECT 15.540 16.650 17.840 16.830 ;
        RECT 21.050 16.650 21.550 17.000 ;
        RECT 15.540 16.350 21.550 16.650 ;
        RECT 31.900 19.050 32.400 20.800 ;
        RECT 73.400 19.050 73.900 24.400 ;
        RECT 31.900 18.550 82.700 19.050 ;
        RECT 31.900 15.800 32.300 18.550 ;
        RECT 37.350 15.800 37.750 18.550 ;
        RECT 42.800 15.800 43.200 18.550 ;
        RECT 52.300 15.800 52.700 18.550 ;
        RECT 61.900 15.800 62.300 18.550 ;
        RECT 67.350 15.800 67.750 18.550 ;
        RECT 72.800 15.800 73.200 18.550 ;
        RECT 82.300 15.800 82.700 18.550 ;
        RECT 92.000 -10.200 92.310 -9.710 ;
        RECT 83.600 -10.220 84.050 -10.200 ;
        RECT 87.700 -10.220 88.150 -10.200 ;
        RECT 91.800 -10.220 92.550 -10.200 ;
        RECT 96.200 -10.220 96.650 -10.200 ;
        RECT 100.300 -10.220 100.750 -10.200 ;
        RECT 79.940 -10.700 104.420 -10.220 ;
        RECT 21.700 -13.850 22.100 -11.600 ;
        RECT 26.000 -13.850 26.400 -11.600 ;
        RECT 28.900 -13.850 29.300 -11.600 ;
        RECT 31.800 -13.850 32.200 -11.600 ;
        RECT 36.100 -13.850 36.500 -11.600 ;
        RECT 40.400 -13.850 40.800 -11.600 ;
        RECT 43.300 -13.850 43.700 -11.600 ;
        RECT 46.200 -13.850 46.600 -11.600 ;
        RECT 50.500 -13.850 50.900 -11.600 ;
        RECT 54.800 -13.850 55.200 -11.600 ;
        RECT 57.700 -13.850 58.100 -11.600 ;
        RECT 60.600 -13.850 61.000 -11.600 ;
        RECT 21.700 -14.250 61.000 -13.850 ;
        RECT 81.950 -14.200 82.350 -13.600 ;
        RECT 99.760 -14.100 100.235 -10.700 ;
        RECT 99.650 -14.200 100.350 -14.100 ;
        RECT 81.750 -14.220 83.750 -14.200 ;
        RECT 91.100 -14.220 93.000 -14.200 ;
        RECT 94.350 -14.220 95.650 -14.200 ;
        RECT 96.950 -14.220 100.350 -14.200 ;
        RECT -16.950 -15.280 -16.400 -15.250 ;
        RECT -15.800 -15.280 -15.400 -14.780 ;
        RECT -16.950 -15.300 -15.100 -15.280 ;
        RECT -16.950 -15.780 -13.370 -15.300 ;
        RECT -11.770 -15.780 -2.110 -15.300 ;
        RECT -0.300 -15.780 1.540 -15.300 ;
        RECT -16.950 -15.800 -16.400 -15.780 ;
        RECT -15.750 -20.480 -15.350 -19.980 ;
        RECT -15.750 -20.510 -15.050 -20.480 ;
        RECT -15.750 -20.990 -13.680 -20.510 ;
        RECT -9.500 -20.830 -9.150 -15.780 ;
        RECT 39.650 -16.050 40.050 -14.250 ;
        RECT 60.600 -16.050 61.000 -14.250 ;
        RECT 79.940 -14.700 100.350 -14.220 ;
        RECT 99.650 -14.800 100.350 -14.700 ;
        RECT 39.650 -16.450 64.550 -16.050 ;
        RECT 28.990 -17.870 29.300 -17.370 ;
        RECT 29.540 -18.300 31.840 -17.820 ;
        RECT 39.650 -18.700 40.050 -16.450 ;
        RECT 42.550 -18.700 42.950 -16.450 ;
        RECT 45.450 -18.700 45.850 -16.450 ;
        RECT 49.750 -18.700 50.150 -16.450 ;
        RECT 54.050 -18.700 54.450 -16.450 ;
        RECT 56.950 -18.700 57.350 -16.450 ;
        RECT 59.850 -18.700 60.250 -16.450 ;
        RECT 64.150 -18.700 64.550 -16.450 ;
        RECT -3.400 -20.980 -2.900 -20.580 ;
        RECT -15.750 -21.030 -15.050 -20.990 ;
        RECT -7.050 -21.460 -0.630 -20.980 ;
        RECT -3.850 -21.480 -2.450 -21.460 ;
        RECT -14.200 -23.430 -12.820 -22.950 ;
        RECT -11.730 -23.430 -2.070 -22.950 ;
        RECT -0.140 -23.430 1.700 -22.950 ;
        RECT -1.000 -23.830 -0.500 -23.430 ;
        RECT 28.950 -29.550 44.450 -29.050 ;
        RECT 43.950 -33.000 44.450 -29.550 ;
        RECT 49.250 -30.750 49.550 -30.250 ;
        RECT 47.140 -31.300 48.980 -30.820 ;
        RECT 43.950 -33.500 50.800 -33.000 ;
        RECT 52.950 -33.500 53.350 -33.000 ;
        RECT 50.300 -37.400 50.800 -33.500 ;
        RECT 54.890 -33.650 57.190 -33.520 ;
        RECT 59.490 -33.600 66.850 -33.520 ;
        RECT 59.490 -33.650 70.150 -33.600 ;
        RECT 54.890 -34.000 70.150 -33.650 ;
        RECT 50.300 -37.900 52.350 -37.400 ;
        RECT 52.690 -38.200 55.450 -37.720 ;
        RECT 58.090 -37.750 67.750 -37.720 ;
        RECT 69.700 -37.750 70.150 -34.000 ;
        RECT 58.090 -38.200 70.150 -37.750 ;
        RECT 77.550 -37.330 77.950 -36.830 ;
        RECT 77.550 -37.350 78.250 -37.330 ;
        RECT 77.550 -37.830 79.980 -37.350 ;
        RECT 81.580 -37.830 91.240 -37.350 ;
        RECT 93.050 -37.830 94.890 -37.350 ;
        RECT 18.100 -43.800 18.580 -41.990 ;
        RECT 18.100 -44.150 18.600 -43.800 ;
        RECT 29.850 -43.900 30.250 -39.900 ;
        RECT 36.900 -43.900 37.300 -41.500 ;
        RECT 77.600 -42.530 78.000 -42.030 ;
        RECT 77.600 -42.560 78.300 -42.530 ;
        RECT 77.600 -43.040 79.670 -42.560 ;
        RECT 83.850 -42.880 84.200 -37.830 ;
        RECT 89.950 -43.030 90.450 -42.630 ;
        RECT 77.600 -43.080 78.300 -43.040 ;
        RECT 86.300 -43.510 92.720 -43.030 ;
        RECT 89.500 -43.530 90.900 -43.510 ;
        RECT 18.100 -44.550 19.100 -44.150 ;
        RECT 29.850 -44.300 37.300 -43.900 ;
        RECT 18.100 -45.300 18.600 -44.550 ;
        RECT 18.100 -46.670 18.580 -45.300 ;
        RECT 17.100 -49.850 17.750 -49.750 ;
        RECT 18.150 -49.850 18.550 -46.670 ;
        RECT 25.400 -49.850 25.800 -47.450 ;
        RECT 29.850 -47.850 30.250 -44.300 ;
        RECT 50.300 -49.100 50.800 -44.700 ;
        RECT 52.950 -45.200 53.350 -44.700 ;
        RECT 79.150 -45.000 79.650 -44.500 ;
        RECT 54.890 -45.350 57.190 -45.220 ;
        RECT 59.490 -45.300 66.850 -45.220 ;
        RECT 59.490 -45.350 70.150 -45.300 ;
        RECT 54.890 -45.700 70.150 -45.350 ;
        RECT 79.150 -45.480 80.530 -45.000 ;
        RECT 81.620 -45.480 91.280 -45.000 ;
        RECT 93.210 -45.480 95.050 -45.000 ;
        RECT 38.515 -49.470 40.620 -49.220 ;
        RECT 50.300 -49.600 52.350 -49.100 ;
        RECT 17.100 -50.250 27.600 -49.850 ;
        RECT 52.690 -49.900 55.450 -49.420 ;
        RECT 58.090 -49.450 67.750 -49.420 ;
        RECT 69.700 -49.450 70.150 -45.700 ;
        RECT 92.350 -45.880 92.850 -45.480 ;
        RECT 58.090 -49.900 70.150 -49.450 ;
        RECT 17.100 -50.400 17.750 -50.250 ;
        RECT 48.550 -55.650 50.200 -54.650 ;
      LAYER met2 ;
        RECT -24.850 24.400 -6.400 24.900 ;
        RECT -24.850 -15.250 -24.350 24.400 ;
        RECT 99.650 -14.800 100.350 -14.100 ;
        RECT -26.425 -15.800 -16.400 -15.250 ;
        RECT -24.850 -49.750 -24.350 -15.800 ;
        RECT 75.600 -44.500 79.650 -44.000 ;
        RECT -24.850 -50.400 17.750 -49.750 ;
        RECT 48.550 -55.000 50.200 -54.650 ;
        RECT 75.600 -55.000 76.100 -44.500 ;
        RECT 79.150 -45.000 79.650 -44.500 ;
        RECT 99.650 -55.000 100.150 -14.800 ;
        RECT 48.550 -55.500 100.150 -55.000 ;
        RECT 48.550 -55.650 50.200 -55.500 ;
    END
  END GND
  PIN Vbs_12
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 26.000 -32.350 26.300 -31.850 ;
        RECT 40.550 -32.400 41.050 -31.900 ;
      LAYER met1 ;
        RECT 15.650 -29.500 26.300 -29.000 ;
        RECT 25.800 -29.900 26.300 -29.500 ;
        RECT 25.800 -30.400 41.050 -29.900 ;
        RECT 25.800 -32.350 26.300 -30.400 ;
        RECT 40.550 -32.400 41.050 -30.400 ;
    END
  END Vbs_12
  PIN VCCA
    ANTENNADIFFAREA 66.559998 ;
    PORT
      LAYER nwell ;
        RECT -7.100 31.850 82.900 37.650 ;
        RECT 22.900 5.800 82.900 11.600 ;
        RECT 24.500 -34.950 26.900 -32.350 ;
        RECT 28.250 -34.950 32.450 -32.350 ;
      LAYER li1 ;
        RECT -6.200 38.150 89.550 38.550 ;
        RECT -6.900 36.800 -6.500 37.300 ;
        RECT -6.200 32.250 -5.800 38.150 ;
        RECT 1.900 32.250 2.300 38.150 ;
        RECT 2.600 36.800 3.000 37.300 ;
        RECT 3.300 32.250 3.700 38.150 ;
        RECT 8.050 36.800 8.450 37.300 ;
        RECT 8.750 32.250 9.150 38.150 ;
        RECT 13.500 36.800 13.900 37.300 ;
        RECT 14.200 32.250 14.600 38.150 ;
        RECT 22.300 32.250 22.700 38.150 ;
        RECT 23.100 36.800 23.500 37.300 ;
        RECT 23.800 32.250 24.200 38.150 ;
        RECT 31.900 32.250 32.300 38.150 ;
        RECT 32.600 36.800 33.000 37.300 ;
        RECT 33.300 32.250 33.700 38.150 ;
        RECT 38.050 36.800 38.450 37.300 ;
        RECT 38.750 32.250 39.150 38.150 ;
        RECT 43.500 36.800 43.900 37.300 ;
        RECT 44.200 32.250 44.600 38.150 ;
        RECT 52.300 32.250 52.700 38.150 ;
        RECT 53.100 36.800 53.500 37.300 ;
        RECT 53.800 32.250 54.200 38.150 ;
        RECT 61.900 32.250 62.300 38.150 ;
        RECT 62.600 36.800 63.000 37.300 ;
        RECT 63.300 32.250 63.700 38.150 ;
        RECT 68.050 36.800 68.450 37.300 ;
        RECT 68.750 32.250 69.150 38.150 ;
        RECT 73.500 36.800 73.900 37.300 ;
        RECT 74.200 32.250 74.600 38.150 ;
        RECT 82.300 32.250 82.700 38.150 ;
        RECT 23.100 5.300 23.500 11.200 ;
        RECT 31.200 5.300 31.600 11.200 ;
        RECT 31.900 6.150 32.300 6.650 ;
        RECT 36.650 5.300 37.050 11.200 ;
        RECT 37.350 6.150 37.750 6.650 ;
        RECT 42.100 5.300 42.500 11.200 ;
        RECT 42.800 6.150 43.200 6.650 ;
        RECT 43.500 5.300 43.900 11.200 ;
        RECT 51.600 5.300 52.000 11.200 ;
        RECT 52.300 6.150 52.700 6.650 ;
        RECT 53.100 5.300 53.500 11.200 ;
        RECT 61.200 5.300 61.600 11.200 ;
        RECT 61.900 6.150 62.300 6.650 ;
        RECT 66.650 5.300 67.050 11.200 ;
        RECT 67.350 6.150 67.750 6.650 ;
        RECT 72.100 5.300 72.500 11.200 ;
        RECT 72.800 6.150 73.200 6.650 ;
        RECT 73.500 5.300 73.900 11.200 ;
        RECT 81.600 5.300 82.000 11.200 ;
        RECT 82.300 6.150 82.700 6.650 ;
        RECT 88.450 5.300 88.950 38.150 ;
        RECT 23.100 4.900 88.950 5.300 ;
        RECT 13.500 -31.250 31.350 -30.850 ;
        RECT 24.700 -33.250 25.100 -31.250 ;
        RECT 25.400 -34.550 25.800 -31.250 ;
        RECT 28.450 -33.200 28.850 -31.250 ;
        RECT 29.150 -34.550 29.550 -32.750 ;
        RECT 30.950 -34.550 31.350 -31.250 ;
      LAYER met1 ;
        RECT -10.400 39.550 89.550 40.050 ;
        RECT -6.900 36.800 -6.500 39.550 ;
        RECT 2.600 36.800 3.000 39.550 ;
        RECT 8.050 36.800 8.450 39.550 ;
        RECT 13.500 36.800 13.900 39.550 ;
        RECT 23.100 36.800 23.500 39.550 ;
        RECT 32.600 36.800 33.000 39.550 ;
        RECT 38.050 36.800 38.450 39.550 ;
        RECT 43.500 36.800 43.900 39.550 ;
        RECT 53.100 36.800 53.500 39.550 ;
        RECT 62.600 36.800 63.000 39.550 ;
        RECT 68.050 36.800 68.450 39.550 ;
        RECT 73.500 36.800 73.900 39.550 ;
        RECT 31.900 3.900 32.300 6.650 ;
        RECT 37.350 3.900 37.750 6.650 ;
        RECT 42.800 3.900 43.200 6.650 ;
        RECT 52.300 3.900 52.700 6.650 ;
        RECT 61.900 3.900 62.300 6.650 ;
        RECT 67.350 3.900 67.750 6.650 ;
        RECT 72.800 3.900 73.200 6.650 ;
        RECT 82.300 3.900 82.700 6.650 ;
        RECT 86.950 3.900 87.450 39.550 ;
        RECT 31.900 3.400 87.450 3.900 ;
        RECT 31.900 -0.300 32.300 3.400 ;
        RECT 13.500 -0.700 32.300 -0.300 ;
        RECT 13.500 -31.250 13.900 -0.700 ;
        RECT 24.700 -33.250 25.100 -32.750 ;
        RECT 28.450 -33.200 28.850 -32.700 ;
        RECT 29.150 -32.900 29.550 -32.750 ;
        RECT 30.950 -32.900 31.350 -32.750 ;
        RECT 29.150 -33.400 31.350 -32.900 ;
        RECT 29.150 -33.550 29.550 -33.400 ;
        RECT 30.950 -33.550 31.350 -33.400 ;
    END
  END VCCA
  PIN Vbs_34
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER li1 ;
        RECT 29.750 -32.350 30.750 -31.850 ;
        RECT 35.050 -32.350 37.350 -31.850 ;
      LAYER met1 ;
        RECT 32.900 -31.850 33.400 -30.950 ;
        RECT 29.550 -32.350 37.350 -31.850 ;
    END
  END Vbs_34
  OBS
      LAYER nwell ;
        RECT 21.500 -9.350 64.700 -5.550 ;
        RECT 35.950 -24.750 64.750 -20.950 ;
        RECT 33.750 -34.950 37.950 -32.350 ;
        RECT 39.250 -35.000 41.650 -32.400 ;
      LAYER pwell ;
        RECT 67.750 -37.900 69.400 -36.950 ;
      LAYER nwell ;
        RECT 24.850 -44.200 28.150 -39.400 ;
        RECT 38.700 -44.250 42.000 -39.450 ;
      LAYER pwell ;
        RECT 67.750 -49.600 69.400 -48.650 ;
      LAYER li1 ;
        RECT -5.000 31.400 -3.800 32.050 ;
        RECT -6.200 26.300 -5.800 31.200 ;
        RECT -2.150 30.850 -1.750 37.250 ;
        RECT -1.300 31.400 -0.100 32.050 ;
        RECT 4.850 31.950 6.050 32.050 ;
        RECT 0.700 31.450 6.050 31.950 ;
        RECT 0.700 30.850 1.200 31.450 ;
        RECT 4.850 31.400 6.050 31.450 ;
        RECT 7.350 32.000 7.750 37.250 ;
        RECT 9.700 32.000 10.900 32.050 ;
        RECT 7.350 31.500 10.900 32.000 ;
        RECT -2.150 30.350 1.200 30.850 ;
        RECT -2.150 27.200 -1.750 30.350 ;
        RECT 1.900 26.300 2.300 31.200 ;
        RECT 3.300 26.300 3.700 31.200 ;
        RECT 7.350 27.200 7.750 31.500 ;
        RECT 9.700 31.400 10.900 31.500 ;
        RECT 8.750 26.300 9.150 31.200 ;
        RECT 12.800 27.200 13.200 37.250 ;
        RECT 15.400 31.400 16.600 32.050 ;
        RECT 14.200 26.300 14.600 31.200 ;
        RECT 18.250 27.200 18.650 37.250 ;
        RECT 19.100 31.400 20.300 32.050 ;
        RECT 25.000 31.400 26.200 32.050 ;
        RECT 22.300 26.300 22.700 31.200 ;
        RECT 23.800 26.300 24.200 31.200 ;
        RECT 27.850 30.850 28.250 37.250 ;
        RECT 28.700 31.400 29.900 32.050 ;
        RECT 34.850 31.950 36.050 32.050 ;
        RECT 30.700 31.450 36.050 31.950 ;
        RECT 30.700 30.850 31.200 31.450 ;
        RECT 34.850 31.400 36.050 31.450 ;
        RECT 37.350 32.000 37.750 37.250 ;
        RECT 39.700 32.000 40.900 32.050 ;
        RECT 37.350 31.500 40.900 32.000 ;
        RECT 27.850 30.350 31.200 30.850 ;
        RECT 27.850 27.200 28.250 30.350 ;
        RECT 31.900 26.300 32.300 31.200 ;
        RECT 33.300 26.300 33.700 31.200 ;
        RECT 37.350 27.200 37.750 31.500 ;
        RECT 39.700 31.400 40.900 31.500 ;
        RECT 38.750 26.300 39.150 31.200 ;
        RECT 42.800 27.200 43.200 37.250 ;
        RECT 45.400 31.400 46.600 32.050 ;
        RECT 44.200 26.300 44.600 31.200 ;
        RECT 48.250 27.200 48.650 37.250 ;
        RECT 49.100 31.400 50.300 32.050 ;
        RECT 55.000 31.400 56.200 32.050 ;
        RECT 52.300 26.300 52.700 31.200 ;
        RECT 53.800 26.300 54.200 31.200 ;
        RECT 57.850 30.850 58.250 37.250 ;
        RECT 58.700 31.400 59.900 32.050 ;
        RECT 64.850 31.950 66.050 32.050 ;
        RECT 60.700 31.450 66.050 31.950 ;
        RECT 60.700 30.850 61.200 31.450 ;
        RECT 64.850 31.400 66.050 31.450 ;
        RECT 67.350 32.000 67.750 37.250 ;
        RECT 69.700 32.000 70.900 32.050 ;
        RECT 67.350 31.500 70.900 32.000 ;
        RECT 57.850 30.350 61.200 30.850 ;
        RECT 57.850 27.200 58.250 30.350 ;
        RECT 61.900 26.300 62.300 31.200 ;
        RECT 63.300 26.300 63.700 31.200 ;
        RECT 67.350 27.200 67.750 31.500 ;
        RECT 69.700 31.400 70.900 31.500 ;
        RECT 68.750 26.300 69.150 31.200 ;
        RECT 72.800 27.200 73.200 37.250 ;
        RECT 75.400 31.400 76.600 32.050 ;
        RECT 74.200 26.300 74.600 31.200 ;
        RECT 78.250 27.200 78.650 37.250 ;
        RECT 79.100 31.400 80.300 32.050 ;
        RECT 82.300 26.300 82.700 31.200 ;
        RECT -6.200 25.900 82.700 26.300 ;
        RECT 16.850 22.880 17.250 22.900 ;
        RECT 16.700 22.850 17.250 22.880 ;
        RECT 23.850 22.850 24.350 25.900 ;
        RECT 16.700 22.800 24.350 22.850 ;
        RECT 14.885 22.480 24.350 22.800 ;
        RECT 16.700 22.450 24.350 22.480 ;
        RECT 16.700 22.400 17.250 22.450 ;
        RECT 23.850 21.400 24.350 22.450 ;
        RECT 23.850 21.330 25.100 21.400 ;
        RECT 23.850 21.250 25.200 21.330 ;
        RECT 23.850 20.930 27.015 21.250 ;
        RECT 23.850 20.850 25.200 20.930 ;
        RECT 23.850 20.800 25.100 20.850 ;
        RECT 15.625 18.655 15.885 19.055 ;
        RECT 17.160 18.715 17.755 19.055 ;
        RECT 15.625 18.485 16.990 18.655 ;
        RECT 16.255 17.415 16.990 18.485 ;
        RECT 15.625 17.245 16.990 17.415 ;
        RECT 17.160 17.395 17.335 18.715 ;
        RECT 23.850 17.550 24.350 20.800 ;
        RECT 81.500 17.550 82.000 25.900 ;
        RECT 15.625 16.845 15.885 17.245 ;
        RECT 17.160 16.845 17.755 17.395 ;
        RECT 23.100 17.150 82.000 17.550 ;
        RECT 23.100 12.250 23.500 17.150 ;
        RECT 25.500 11.400 26.700 12.050 ;
        RECT 27.150 6.200 27.550 16.250 ;
        RECT 31.200 12.250 31.600 17.150 ;
        RECT 29.200 11.400 30.400 12.050 ;
        RECT 32.600 6.200 33.000 16.250 ;
        RECT 36.650 12.250 37.050 17.150 ;
        RECT 34.900 11.950 36.100 12.050 ;
        RECT 38.050 11.950 38.450 16.250 ;
        RECT 42.100 12.250 42.500 17.150 ;
        RECT 43.500 12.250 43.900 17.150 ;
        RECT 47.550 13.100 47.950 16.250 ;
        RECT 44.600 12.600 47.950 13.100 ;
        RECT 34.900 11.450 38.450 11.950 ;
        RECT 34.900 11.400 36.100 11.450 ;
        RECT 38.050 6.200 38.450 11.450 ;
        RECT 39.750 12.000 40.950 12.050 ;
        RECT 44.600 12.000 45.100 12.600 ;
        RECT 39.750 11.500 45.100 12.000 ;
        RECT 39.750 11.400 40.950 11.500 ;
        RECT 45.900 11.400 47.100 12.050 ;
        RECT 47.550 6.200 47.950 12.600 ;
        RECT 51.600 12.250 52.000 17.150 ;
        RECT 53.100 12.250 53.500 17.150 ;
        RECT 49.600 11.400 50.800 12.050 ;
        RECT 55.500 11.400 56.700 12.050 ;
        RECT 57.150 6.200 57.550 16.250 ;
        RECT 61.200 12.250 61.600 17.150 ;
        RECT 59.200 11.400 60.400 12.050 ;
        RECT 62.600 6.200 63.000 16.250 ;
        RECT 66.650 12.250 67.050 17.150 ;
        RECT 64.900 11.950 66.100 12.050 ;
        RECT 68.050 11.950 68.450 16.250 ;
        RECT 72.100 12.250 72.500 17.150 ;
        RECT 73.500 12.250 73.900 17.150 ;
        RECT 77.550 13.100 77.950 16.250 ;
        RECT 74.600 12.600 77.950 13.100 ;
        RECT 64.900 11.450 68.450 11.950 ;
        RECT 64.900 11.400 66.100 11.450 ;
        RECT 68.050 6.200 68.450 11.450 ;
        RECT 69.750 12.000 70.950 12.050 ;
        RECT 74.600 12.000 75.100 12.600 ;
        RECT 69.750 11.500 75.100 12.000 ;
        RECT 69.750 11.400 70.950 11.500 ;
        RECT 75.900 11.400 77.100 12.050 ;
        RECT 77.550 6.200 77.950 12.600 ;
        RECT 81.600 12.250 82.000 17.150 ;
        RECT 79.600 11.400 80.800 12.050 ;
        RECT 22.400 -5.050 66.300 -4.650 ;
        RECT 21.700 -6.400 22.100 -5.900 ;
        RECT 22.400 -8.950 22.800 -5.050 ;
        RECT 23.050 -9.750 23.500 -9.300 ;
        RECT 23.800 -12.050 24.200 -5.950 ;
        RECT 25.200 -8.950 25.600 -5.050 ;
        RECT 26.000 -6.500 26.400 -6.000 ;
        RECT 26.700 -8.950 27.100 -5.050 ;
        RECT 28.100 -9.300 28.500 -5.950 ;
        RECT 28.900 -6.500 29.300 -6.000 ;
        RECT 29.600 -8.950 30.000 -5.050 ;
        RECT 24.450 -9.750 24.900 -9.300 ;
        RECT 27.350 -9.700 27.750 -9.300 ;
        RECT 28.100 -9.700 30.650 -9.300 ;
        RECT 28.100 -12.050 28.500 -9.700 ;
        RECT 31.000 -12.050 31.400 -5.950 ;
        RECT 31.800 -6.400 32.200 -5.900 ;
        RECT 32.500 -8.950 32.900 -5.050 ;
        RECT 33.150 -9.750 33.600 -9.300 ;
        RECT 33.900 -12.050 34.300 -5.950 ;
        RECT 35.300 -8.950 35.700 -5.050 ;
        RECT 36.100 -6.400 36.500 -5.900 ;
        RECT 36.800 -8.950 37.200 -5.050 ;
        RECT 34.550 -9.750 35.000 -9.300 ;
        RECT 37.450 -9.750 37.900 -9.300 ;
        RECT 38.200 -12.050 38.600 -5.950 ;
        RECT 39.600 -8.950 40.000 -5.050 ;
        RECT 40.400 -6.500 40.800 -6.000 ;
        RECT 41.100 -8.950 41.500 -5.050 ;
        RECT 42.500 -9.300 42.900 -5.950 ;
        RECT 43.300 -6.500 43.700 -6.000 ;
        RECT 44.000 -8.950 44.400 -5.050 ;
        RECT 38.850 -9.750 39.300 -9.300 ;
        RECT 41.750 -9.700 42.150 -9.300 ;
        RECT 42.500 -9.700 45.050 -9.300 ;
        RECT 42.500 -12.050 42.900 -9.700 ;
        RECT 45.400 -12.050 45.800 -5.950 ;
        RECT 46.200 -6.400 46.600 -5.900 ;
        RECT 46.900 -8.950 47.300 -5.050 ;
        RECT 47.550 -9.750 48.000 -9.300 ;
        RECT 48.300 -12.050 48.700 -5.950 ;
        RECT 49.700 -8.950 50.100 -5.050 ;
        RECT 50.500 -6.400 50.900 -5.900 ;
        RECT 51.200 -8.950 51.600 -5.050 ;
        RECT 48.950 -9.750 49.400 -9.300 ;
        RECT 51.850 -9.750 52.300 -9.300 ;
        RECT 52.600 -12.050 53.000 -5.950 ;
        RECT 54.000 -8.950 54.400 -5.050 ;
        RECT 54.800 -6.500 55.200 -6.000 ;
        RECT 55.500 -8.950 55.900 -5.050 ;
        RECT 56.900 -9.300 57.300 -5.950 ;
        RECT 57.700 -6.500 58.100 -6.000 ;
        RECT 58.400 -8.950 58.800 -5.050 ;
        RECT 53.250 -9.750 53.700 -9.300 ;
        RECT 56.150 -9.700 56.550 -9.300 ;
        RECT 56.900 -9.700 59.450 -9.300 ;
        RECT 56.900 -12.050 57.300 -9.700 ;
        RECT 59.800 -12.050 60.200 -5.950 ;
        RECT 60.600 -6.400 61.000 -5.900 ;
        RECT 61.300 -8.950 61.700 -5.050 ;
        RECT 61.950 -9.750 62.400 -9.300 ;
        RECT 62.700 -12.050 63.100 -5.950 ;
        RECT 64.100 -8.950 64.500 -5.050 ;
        RECT 63.350 -9.750 63.800 -9.300 ;
        RECT -15.035 -13.835 -14.865 -13.075 ;
        RECT -15.035 -14.005 -14.320 -13.835 ;
        RECT -14.150 -13.980 -13.895 -13.075 ;
        RECT -11.595 -13.575 -11.425 -13.075 ;
        RECT -11.595 -13.745 -10.930 -13.575 ;
        RECT -16.500 -14.180 -16.000 -14.150 ;
        RECT -16.500 -14.530 -14.750 -14.180 ;
        RECT -14.490 -14.215 -14.320 -14.005 ;
        RECT -16.500 -14.600 -16.000 -14.530 ;
        RECT -15.125 -14.555 -14.770 -14.530 ;
        RECT -14.490 -14.545 -14.235 -14.215 ;
        RECT -14.065 -14.230 -13.895 -13.980 ;
        RECT -11.680 -14.230 -11.330 -13.915 ;
        RECT -14.065 -14.430 -11.330 -14.230 ;
        RECT -14.490 -14.735 -14.320 -14.545 ;
        RECT -14.065 -14.710 -13.895 -14.430 ;
        RECT -11.680 -14.565 -11.330 -14.430 ;
        RECT -15.035 -14.905 -14.320 -14.735 ;
        RECT -15.035 -15.285 -14.865 -14.905 ;
        RECT -14.150 -15.285 -13.895 -14.710 ;
        RECT -11.160 -14.735 -10.930 -13.745 ;
        RECT -11.595 -14.905 -10.930 -14.735 ;
        RECT -11.595 -15.195 -11.425 -14.905 ;
        RECT -10.755 -15.195 -10.530 -13.075 ;
        RECT -9.815 -13.575 -9.645 -13.075 ;
        RECT -9.410 -13.290 -8.580 -13.120 ;
        RECT -10.340 -13.745 -9.645 -13.575 ;
        RECT -10.340 -14.715 -10.170 -13.745 ;
        RECT -10.000 -14.535 -9.590 -13.915 ;
        RECT -9.420 -13.965 -8.920 -13.585 ;
        RECT -10.340 -14.905 -9.645 -14.715 ;
        RECT -9.420 -14.835 -9.200 -13.965 ;
        RECT -8.750 -14.135 -8.580 -13.290 ;
        RECT -7.780 -13.455 -7.610 -13.165 ;
        RECT -6.640 -13.375 -6.010 -13.125 ;
        RECT -6.180 -13.455 -6.010 -13.375 ;
        RECT -5.210 -13.455 -4.970 -13.165 ;
        RECT -8.410 -13.705 -7.040 -13.455 ;
        RECT -8.410 -13.965 -8.160 -13.705 ;
        RECT -7.650 -14.135 -7.400 -13.975 ;
        RECT -8.750 -14.305 -7.400 -14.135 ;
        RECT -8.750 -14.345 -8.330 -14.305 ;
        RECT -9.020 -14.895 -8.670 -14.525 ;
        RECT -9.815 -15.235 -9.645 -14.905 ;
        RECT -8.500 -15.075 -8.330 -14.345 ;
        RECT -7.230 -14.475 -7.040 -13.705 ;
        RECT -8.160 -14.805 -7.750 -14.475 ;
        RECT -9.345 -15.275 -8.330 -15.075 ;
        RECT -7.460 -14.815 -7.040 -14.475 ;
        RECT -6.870 -13.885 -6.350 -13.575 ;
        RECT -6.180 -13.625 -4.970 -13.455 ;
        RECT -6.870 -14.645 -6.700 -13.885 ;
        RECT -6.530 -14.475 -6.350 -14.065 ;
        RECT -6.180 -14.135 -6.010 -13.625 ;
        RECT -4.240 -13.775 -4.070 -13.165 ;
        RECT -3.800 -13.625 -3.470 -13.115 ;
        RECT -4.240 -13.795 -3.920 -13.775 ;
        RECT -5.840 -13.965 -3.920 -13.795 ;
        RECT -6.180 -14.305 -4.280 -14.135 ;
        RECT -5.950 -14.645 -5.620 -14.525 ;
        RECT -6.870 -14.815 -5.620 -14.645 ;
        RECT -7.460 -15.245 -7.210 -14.815 ;
        RECT -5.450 -15.065 -5.280 -14.305 ;
        RECT -4.610 -14.365 -4.280 -14.305 ;
        RECT -5.090 -14.535 -4.760 -14.475 ;
        RECT -5.090 -14.805 -4.430 -14.535 ;
        RECT -4.110 -14.860 -3.920 -13.965 ;
        RECT -6.130 -15.235 -5.280 -15.065 ;
        RECT -4.240 -15.190 -3.920 -14.860 ;
        RECT -3.720 -14.215 -3.470 -13.625 ;
        RECT -2.825 -13.885 -2.570 -13.215 ;
        RECT -2.750 -14.180 -2.570 -13.885 ;
        RECT -0.125 -13.835 0.045 -13.075 ;
        RECT -0.125 -14.005 0.590 -13.835 ;
        RECT 0.760 -13.980 1.015 -13.075 ;
        RECT -2.750 -14.185 -0.200 -14.180 ;
        RECT -3.720 -14.545 -2.920 -14.215 ;
        RECT -3.720 -15.195 -3.470 -14.545 ;
        RECT -2.750 -14.555 0.140 -14.185 ;
        RECT 0.420 -14.215 0.590 -14.005 ;
        RECT 0.420 -14.545 0.675 -14.215 ;
        RECT -2.750 -14.580 -0.200 -14.555 ;
        RECT -2.750 -14.745 -2.570 -14.580 ;
        RECT 0.420 -14.735 0.590 -14.545 ;
        RECT 0.845 -14.710 1.015 -13.980 ;
        RECT -2.825 -15.275 -2.570 -14.745 ;
        RECT -0.125 -14.905 0.590 -14.735 ;
        RECT -0.125 -15.285 0.045 -14.905 ;
        RECT 0.760 -15.285 1.015 -14.710 ;
        RECT 29.625 -15.995 29.885 -15.595 ;
        RECT 31.160 -15.600 31.755 -15.595 ;
        RECT 31.160 -15.900 34.050 -15.600 ;
        RECT 31.160 -15.935 31.755 -15.900 ;
        RECT 29.625 -16.165 30.990 -15.995 ;
        RECT 30.255 -17.235 30.990 -16.165 ;
        RECT 29.625 -17.405 30.990 -17.235 ;
        RECT 31.160 -17.255 31.335 -15.935 ;
        RECT 29.625 -17.805 29.885 -17.405 ;
        RECT 31.160 -17.805 31.755 -17.255 ;
        RECT -14.535 -19.265 -14.205 -18.285 ;
        RECT -14.455 -19.480 -14.205 -19.265 ;
        RECT -6.965 -19.435 -6.585 -18.755 ;
        RECT -5.655 -19.265 -5.325 -18.755 ;
        RECT -4.815 -19.265 -4.415 -18.755 ;
        RECT -5.655 -19.435 -4.415 -19.265 ;
        RECT -14.455 -19.650 -14.200 -19.480 ;
        RECT -14.455 -19.865 -14.205 -19.650 ;
        RECT -14.535 -20.495 -14.205 -19.865 ;
        RECT -6.965 -20.395 -6.795 -19.435 ;
        RECT -6.625 -19.775 -5.320 -19.605 ;
        RECT -4.235 -19.685 -3.915 -18.755 ;
        RECT -2.295 -19.515 -2.125 -18.755 ;
        RECT -2.295 -19.685 -1.580 -19.515 ;
        RECT -1.410 -19.660 -1.155 -18.755 ;
        RECT 33.750 -19.050 34.050 -15.900 ;
        RECT 33.700 -19.450 34.100 -19.050 ;
        RECT -6.625 -20.225 -6.380 -19.775 ;
        RECT -6.210 -20.145 -5.660 -19.945 ;
        RECT -5.490 -19.975 -5.320 -19.775 ;
        RECT -4.545 -19.830 -3.915 -19.685 ;
        RECT -4.545 -19.880 -2.700 -19.830 ;
        RECT -2.385 -19.880 -2.030 -19.865 ;
        RECT -5.490 -20.145 -5.115 -19.975 ;
        RECT -4.945 -20.395 -4.715 -19.895 ;
        RECT -6.965 -20.565 -4.715 -20.395 ;
        RECT -4.545 -20.080 -2.030 -19.880 ;
        RECT -6.415 -20.885 -6.245 -20.565 ;
        RECT -4.545 -20.735 -4.375 -20.080 ;
        RECT -2.385 -20.235 -2.030 -20.080 ;
        RECT -1.750 -19.895 -1.580 -19.685 ;
        RECT -1.750 -20.225 -1.495 -19.895 ;
        RECT -1.750 -20.415 -1.580 -20.225 ;
        RECT -1.325 -20.390 -1.155 -19.660 ;
        RECT -5.330 -20.905 -4.375 -20.735 ;
        RECT -2.295 -20.585 -1.580 -20.415 ;
        RECT -2.295 -20.965 -2.125 -20.585 ;
        RECT -1.410 -20.965 -1.155 -20.390 ;
        RECT 36.850 -21.000 37.300 -20.550 ;
        RECT -13.675 -24.075 -13.345 -23.445 ;
        RECT -11.270 -23.985 -11.015 -23.455 ;
        RECT -13.675 -24.675 -13.425 -24.075 ;
        RECT -13.255 -24.270 -12.925 -24.265 ;
        RECT -11.270 -24.270 -11.090 -23.985 ;
        RECT -10.370 -24.185 -10.120 -23.535 ;
        RECT -13.255 -24.510 -11.090 -24.270 ;
        RECT -13.255 -24.515 -12.925 -24.510 ;
        RECT -13.675 -25.655 -13.345 -24.675 ;
        RECT -11.270 -24.845 -11.090 -24.510 ;
        RECT -10.920 -24.515 -10.120 -24.185 ;
        RECT -11.270 -25.515 -11.015 -24.845 ;
        RECT -10.370 -25.105 -10.120 -24.515 ;
        RECT -9.920 -23.870 -9.600 -23.540 ;
        RECT -8.560 -23.665 -7.710 -23.495 ;
        RECT -9.920 -24.765 -9.730 -23.870 ;
        RECT -9.410 -24.195 -8.750 -23.925 ;
        RECT -9.080 -24.255 -8.750 -24.195 ;
        RECT -9.560 -24.425 -9.230 -24.365 ;
        RECT -8.560 -24.425 -8.390 -23.665 ;
        RECT -6.630 -23.915 -6.380 -23.485 ;
        RECT -8.220 -24.085 -6.970 -23.915 ;
        RECT -8.220 -24.205 -7.890 -24.085 ;
        RECT -9.560 -24.595 -7.660 -24.425 ;
        RECT -9.920 -24.935 -8.000 -24.765 ;
        RECT -9.920 -24.955 -9.600 -24.935 ;
        RECT -10.370 -25.615 -10.040 -25.105 ;
        RECT -9.770 -25.565 -9.600 -24.955 ;
        RECT -7.830 -25.105 -7.660 -24.595 ;
        RECT -7.490 -24.665 -7.310 -24.255 ;
        RECT -7.140 -24.845 -6.970 -24.085 ;
        RECT -8.870 -25.275 -7.660 -25.105 ;
        RECT -7.490 -25.155 -6.970 -24.845 ;
        RECT -6.800 -24.255 -6.380 -23.915 ;
        RECT -5.510 -23.655 -4.495 -23.455 ;
        RECT -6.090 -24.255 -5.680 -23.925 ;
        RECT -6.800 -25.025 -6.610 -24.255 ;
        RECT -5.510 -24.385 -5.340 -23.655 ;
        RECT -4.195 -23.825 -4.025 -23.495 ;
        RECT -5.170 -24.205 -4.820 -23.835 ;
        RECT -5.510 -24.425 -5.090 -24.385 ;
        RECT -6.440 -24.595 -5.090 -24.425 ;
        RECT -6.440 -24.755 -6.190 -24.595 ;
        RECT -5.680 -25.025 -5.430 -24.765 ;
        RECT -6.800 -25.275 -5.430 -25.025 ;
        RECT -8.870 -25.565 -8.630 -25.275 ;
        RECT -7.830 -25.355 -7.660 -25.275 ;
        RECT -7.830 -25.605 -7.200 -25.355 ;
        RECT -6.230 -25.565 -6.060 -25.275 ;
        RECT -5.260 -25.440 -5.090 -24.595 ;
        RECT -4.640 -24.765 -4.420 -23.895 ;
        RECT -4.195 -24.015 -3.500 -23.825 ;
        RECT -4.920 -25.145 -4.420 -24.765 ;
        RECT -4.250 -24.815 -3.840 -24.195 ;
        RECT -3.670 -24.985 -3.500 -24.015 ;
        RECT -4.195 -25.155 -3.500 -24.985 ;
        RECT -5.260 -25.610 -4.430 -25.440 ;
        RECT -4.195 -25.655 -4.025 -25.155 ;
        RECT -3.310 -25.655 -3.085 -23.535 ;
        RECT -2.415 -23.825 -2.245 -23.535 ;
        RECT -2.910 -23.995 -2.245 -23.825 ;
        RECT -2.910 -24.985 -2.680 -23.995 ;
        RECT 0.385 -24.020 0.640 -23.445 ;
        RECT 1.355 -23.825 1.525 -23.445 ;
        RECT 0.810 -23.995 1.525 -23.825 ;
        RECT -2.510 -24.180 -2.160 -24.165 ;
        RECT -2.510 -24.530 -0.600 -24.180 ;
        RECT -2.510 -24.815 -2.160 -24.530 ;
        RECT 0.385 -24.750 0.555 -24.020 ;
        RECT 0.810 -24.185 0.980 -23.995 ;
        RECT 1.950 -24.130 2.850 -24.100 ;
        RECT 1.900 -24.170 2.850 -24.130 ;
        RECT 0.725 -24.515 0.980 -24.185 ;
        RECT 0.810 -24.725 0.980 -24.515 ;
        RECT 1.260 -24.550 2.850 -24.170 ;
        RECT 1.900 -24.580 2.850 -24.550 ;
        RECT 1.950 -24.600 2.850 -24.580 ;
        RECT -2.910 -25.155 -2.245 -24.985 ;
        RECT -2.415 -25.655 -2.245 -25.155 ;
        RECT 0.385 -25.655 0.640 -24.750 ;
        RECT 0.810 -24.895 1.525 -24.725 ;
        RECT 1.355 -25.655 1.525 -24.895 ;
        RECT 36.150 -25.250 36.550 -21.350 ;
        RECT 37.550 -24.350 37.950 -18.250 ;
        RECT 38.250 -21.000 38.700 -20.550 ;
        RECT 38.950 -25.250 39.350 -21.350 ;
        RECT 39.650 -24.400 40.050 -23.900 ;
        RECT 40.450 -24.350 40.850 -18.250 ;
        RECT 43.350 -20.600 43.750 -18.250 ;
        RECT 41.200 -21.000 43.750 -20.600 ;
        RECT 44.100 -21.000 44.500 -20.600 ;
        RECT 46.950 -21.000 47.400 -20.550 ;
        RECT 41.850 -25.250 42.250 -21.350 ;
        RECT 42.550 -24.300 42.950 -23.800 ;
        RECT 43.350 -24.350 43.750 -21.000 ;
        RECT 44.750 -25.250 45.150 -21.350 ;
        RECT 45.450 -24.300 45.850 -23.800 ;
        RECT 46.250 -25.250 46.650 -21.350 ;
        RECT 47.650 -24.350 48.050 -18.250 ;
        RECT 48.350 -21.000 48.800 -20.550 ;
        RECT 51.250 -21.000 51.700 -20.550 ;
        RECT 49.050 -25.250 49.450 -21.350 ;
        RECT 49.750 -24.400 50.150 -23.900 ;
        RECT 50.550 -25.250 50.950 -21.350 ;
        RECT 51.950 -24.350 52.350 -18.250 ;
        RECT 52.650 -21.000 53.100 -20.550 ;
        RECT 53.350 -25.250 53.750 -21.350 ;
        RECT 54.050 -24.400 54.450 -23.900 ;
        RECT 54.850 -24.350 55.250 -18.250 ;
        RECT 57.750 -20.600 58.150 -18.250 ;
        RECT 55.600 -21.000 58.150 -20.600 ;
        RECT 58.500 -21.000 58.900 -20.600 ;
        RECT 61.350 -21.000 61.800 -20.550 ;
        RECT 56.250 -25.250 56.650 -21.350 ;
        RECT 56.950 -24.300 57.350 -23.800 ;
        RECT 57.750 -24.350 58.150 -21.000 ;
        RECT 59.150 -25.250 59.550 -21.350 ;
        RECT 59.850 -24.300 60.250 -23.800 ;
        RECT 60.650 -25.250 61.050 -21.350 ;
        RECT 62.050 -24.350 62.450 -18.250 ;
        RECT 62.750 -21.000 63.200 -20.550 ;
        RECT 63.450 -25.250 63.850 -21.350 ;
        RECT 64.150 -24.400 64.550 -23.900 ;
        RECT 65.900 -25.250 66.300 -5.050 ;
        RECT 80.140 -8.455 80.425 -7.995 ;
        RECT 80.140 -8.675 81.095 -8.455 ;
        RECT 80.885 -9.575 81.095 -8.675 ;
        RECT 80.140 -9.745 81.095 -9.575 ;
        RECT 81.265 -8.845 81.665 -7.995 ;
        RECT 81.855 -8.455 82.135 -7.995 ;
        RECT 81.855 -8.675 82.980 -8.455 ;
        RECT 81.265 -9.405 82.360 -8.845 ;
        RECT 82.530 -9.135 82.980 -8.675 ;
        RECT 83.150 -8.850 83.535 -7.995 ;
        RECT 84.240 -8.455 84.525 -7.995 ;
        RECT 84.240 -8.675 85.195 -8.455 ;
        RECT 84.125 -8.850 84.815 -8.845 ;
        RECT 83.150 -8.965 84.815 -8.850 ;
        RECT 80.140 -10.205 80.425 -9.745 ;
        RECT 81.265 -10.205 81.665 -9.405 ;
        RECT 82.530 -9.465 83.085 -9.135 ;
        RECT 83.255 -9.400 84.815 -8.965 ;
        RECT 82.530 -9.575 82.980 -9.465 ;
        RECT 81.855 -9.745 82.980 -9.575 ;
        RECT 83.255 -9.635 83.535 -9.400 ;
        RECT 84.125 -9.405 84.815 -9.400 ;
        RECT 84.985 -9.575 85.195 -8.675 ;
        RECT 81.855 -10.205 82.135 -9.745 ;
        RECT 83.150 -10.205 83.535 -9.635 ;
        RECT 84.240 -9.745 85.195 -9.575 ;
        RECT 85.365 -8.845 85.765 -7.995 ;
        RECT 85.955 -8.455 86.235 -7.995 ;
        RECT 85.955 -8.675 87.080 -8.455 ;
        RECT 85.365 -9.405 86.460 -8.845 ;
        RECT 86.630 -9.135 87.080 -8.675 ;
        RECT 87.250 -8.850 87.635 -7.995 ;
        RECT 88.340 -8.455 88.625 -7.995 ;
        RECT 88.340 -8.675 89.295 -8.455 ;
        RECT 88.225 -8.850 88.915 -8.845 ;
        RECT 87.250 -8.965 88.915 -8.850 ;
        RECT 84.240 -10.205 84.525 -9.745 ;
        RECT 85.365 -10.205 85.765 -9.405 ;
        RECT 86.630 -9.465 87.185 -9.135 ;
        RECT 87.355 -9.400 88.915 -8.965 ;
        RECT 86.630 -9.575 87.080 -9.465 ;
        RECT 85.955 -9.745 87.080 -9.575 ;
        RECT 87.355 -9.635 87.635 -9.400 ;
        RECT 88.225 -9.405 88.915 -9.400 ;
        RECT 89.085 -9.575 89.295 -8.675 ;
        RECT 85.955 -10.205 86.235 -9.745 ;
        RECT 87.250 -10.205 87.635 -9.635 ;
        RECT 88.340 -9.745 89.295 -9.575 ;
        RECT 89.465 -8.845 89.865 -7.995 ;
        RECT 90.055 -8.455 90.335 -7.995 ;
        RECT 90.055 -8.675 91.180 -8.455 ;
        RECT 89.465 -9.405 90.560 -8.845 ;
        RECT 90.730 -9.135 91.180 -8.675 ;
        RECT 91.350 -8.850 91.735 -7.995 ;
        RECT 92.740 -8.455 93.025 -7.995 ;
        RECT 92.740 -8.675 93.695 -8.455 ;
        RECT 92.625 -8.850 93.315 -8.845 ;
        RECT 91.350 -8.965 93.315 -8.850 ;
        RECT 88.340 -10.205 88.625 -9.745 ;
        RECT 89.465 -10.205 89.865 -9.405 ;
        RECT 90.730 -9.465 91.285 -9.135 ;
        RECT 91.455 -9.400 93.315 -8.965 ;
        RECT 90.730 -9.575 91.180 -9.465 ;
        RECT 90.055 -9.745 91.180 -9.575 ;
        RECT 91.455 -9.635 91.735 -9.400 ;
        RECT 92.625 -9.405 93.315 -9.400 ;
        RECT 93.485 -9.575 93.695 -8.675 ;
        RECT 90.055 -10.205 90.335 -9.745 ;
        RECT 91.350 -10.205 91.735 -9.635 ;
        RECT 92.740 -9.745 93.695 -9.575 ;
        RECT 93.865 -8.845 94.265 -7.995 ;
        RECT 94.455 -8.455 94.735 -7.995 ;
        RECT 94.455 -8.675 95.580 -8.455 ;
        RECT 93.865 -9.405 94.960 -8.845 ;
        RECT 95.130 -9.135 95.580 -8.675 ;
        RECT 95.750 -8.850 96.135 -7.995 ;
        RECT 96.840 -8.455 97.125 -7.995 ;
        RECT 96.840 -8.675 97.795 -8.455 ;
        RECT 96.725 -8.850 97.415 -8.845 ;
        RECT 95.750 -8.965 97.415 -8.850 ;
        RECT 92.740 -10.205 93.025 -9.745 ;
        RECT 93.865 -10.205 94.265 -9.405 ;
        RECT 95.130 -9.465 95.685 -9.135 ;
        RECT 95.855 -9.400 97.415 -8.965 ;
        RECT 95.130 -9.575 95.580 -9.465 ;
        RECT 94.455 -9.745 95.580 -9.575 ;
        RECT 95.855 -9.635 96.135 -9.400 ;
        RECT 96.725 -9.405 97.415 -9.400 ;
        RECT 97.585 -9.575 97.795 -8.675 ;
        RECT 94.455 -10.205 94.735 -9.745 ;
        RECT 95.750 -10.205 96.135 -9.635 ;
        RECT 96.840 -9.745 97.795 -9.575 ;
        RECT 97.965 -8.845 98.365 -7.995 ;
        RECT 98.555 -8.455 98.835 -7.995 ;
        RECT 98.555 -8.675 99.680 -8.455 ;
        RECT 97.965 -9.405 99.060 -8.845 ;
        RECT 99.230 -9.135 99.680 -8.675 ;
        RECT 99.850 -8.850 100.235 -7.995 ;
        RECT 100.940 -8.455 101.225 -7.995 ;
        RECT 100.940 -8.675 101.895 -8.455 ;
        RECT 100.825 -8.850 101.515 -8.845 ;
        RECT 99.850 -8.965 101.515 -8.850 ;
        RECT 96.840 -10.205 97.125 -9.745 ;
        RECT 97.965 -10.205 98.365 -9.405 ;
        RECT 99.230 -9.465 99.785 -9.135 ;
        RECT 99.955 -9.400 101.515 -8.965 ;
        RECT 99.230 -9.575 99.680 -9.465 ;
        RECT 98.555 -9.745 99.680 -9.575 ;
        RECT 99.955 -9.635 100.235 -9.400 ;
        RECT 100.825 -9.405 101.515 -9.400 ;
        RECT 101.685 -9.575 101.895 -8.675 ;
        RECT 98.555 -10.205 98.835 -9.745 ;
        RECT 99.850 -10.205 100.235 -9.635 ;
        RECT 100.940 -9.745 101.895 -9.575 ;
        RECT 102.065 -8.845 102.465 -7.995 ;
        RECT 102.655 -8.455 102.935 -7.995 ;
        RECT 102.655 -8.675 103.780 -8.455 ;
        RECT 102.065 -9.405 103.160 -8.845 ;
        RECT 103.330 -9.135 103.780 -8.675 ;
        RECT 103.950 -8.965 104.335 -7.995 ;
        RECT 100.940 -10.205 101.225 -9.745 ;
        RECT 102.065 -10.205 102.465 -9.405 ;
        RECT 103.330 -9.465 103.885 -9.135 ;
        RECT 103.330 -9.575 103.780 -9.465 ;
        RECT 102.655 -9.745 103.780 -9.575 ;
        RECT 104.055 -9.550 104.335 -8.965 ;
        RECT 104.055 -9.635 105.750 -9.550 ;
        RECT 102.655 -10.205 102.935 -9.745 ;
        RECT 103.950 -9.900 105.750 -9.635 ;
        RECT 103.950 -10.205 104.335 -9.900 ;
        RECT 105.400 -10.900 105.750 -9.900 ;
        RECT 94.800 -11.250 105.750 -10.900 ;
        RECT 80.115 -12.755 80.285 -11.995 ;
        RECT 80.115 -12.925 80.830 -12.755 ;
        RECT 81.000 -12.900 81.255 -11.995 ;
        RECT 83.915 -12.495 84.085 -11.995 ;
        RECT 83.915 -12.665 84.580 -12.495 ;
        RECT 80.025 -13.475 80.380 -13.105 ;
        RECT 80.660 -13.135 80.830 -12.925 ;
        RECT 80.660 -13.465 80.915 -13.135 ;
        RECT 80.660 -13.655 80.830 -13.465 ;
        RECT 81.085 -13.630 81.255 -12.900 ;
        RECT 80.115 -13.825 80.830 -13.655 ;
        RECT 80.115 -14.205 80.285 -13.825 ;
        RECT 81.000 -14.205 81.255 -13.630 ;
        RECT 84.350 -13.655 84.580 -12.665 ;
        RECT 83.915 -13.825 84.580 -13.655 ;
        RECT 83.915 -14.115 84.085 -13.825 ;
        RECT 84.755 -14.115 84.940 -11.995 ;
        RECT 85.615 -12.420 85.865 -11.995 ;
        RECT 86.075 -12.270 87.180 -12.100 ;
        RECT 85.560 -12.550 85.865 -12.420 ;
        RECT 85.110 -13.745 85.390 -12.795 ;
        RECT 85.560 -13.655 85.730 -12.550 ;
        RECT 85.900 -13.335 86.140 -12.740 ;
        RECT 86.310 -12.805 86.840 -12.440 ;
        RECT 86.310 -13.505 86.480 -12.805 ;
        RECT 87.010 -12.885 87.180 -12.270 ;
        RECT 87.690 -12.325 87.940 -11.995 ;
        RECT 88.165 -12.295 89.050 -12.125 ;
        RECT 87.010 -12.975 87.520 -12.885 ;
        RECT 85.560 -13.785 85.785 -13.655 ;
        RECT 85.955 -13.725 86.480 -13.505 ;
        RECT 86.650 -13.145 87.520 -12.975 ;
        RECT 85.615 -13.925 85.785 -13.785 ;
        RECT 86.650 -13.925 86.820 -13.145 ;
        RECT 87.350 -13.215 87.520 -13.145 ;
        RECT 87.030 -13.395 87.230 -13.365 ;
        RECT 87.690 -13.395 87.860 -12.325 ;
        RECT 88.030 -13.215 88.220 -12.495 ;
        RECT 87.030 -13.695 87.860 -13.395 ;
        RECT 88.390 -13.425 88.710 -12.465 ;
        RECT 85.615 -14.095 85.950 -13.925 ;
        RECT 86.145 -14.095 86.820 -13.925 ;
        RECT 87.690 -13.925 87.860 -13.695 ;
        RECT 88.245 -13.755 88.710 -13.425 ;
        RECT 88.880 -13.135 89.050 -12.295 ;
        RECT 89.775 -12.555 90.115 -11.995 ;
        RECT 89.220 -12.930 90.115 -12.555 ;
        RECT 89.925 -13.135 90.115 -12.930 ;
        RECT 93.525 -12.975 93.855 -11.995 ;
        RECT 88.880 -13.465 89.755 -13.135 ;
        RECT 89.925 -13.465 90.675 -13.135 ;
        RECT 88.880 -13.925 89.050 -13.465 ;
        RECT 89.925 -13.635 90.125 -13.465 ;
        RECT 87.690 -14.095 88.095 -13.925 ;
        RECT 88.265 -14.095 89.050 -13.925 ;
        RECT 89.795 -14.160 90.125 -13.635 ;
        RECT 93.590 -13.575 93.760 -12.975 ;
        RECT 93.930 -13.150 94.265 -13.135 ;
        RECT 94.800 -13.150 95.150 -11.250 ;
        RECT 96.165 -12.975 96.495 -11.995 ;
        RECT 97.800 -12.750 108.550 -12.400 ;
        RECT 93.930 -13.385 95.150 -13.150 ;
        RECT 95.745 -13.385 96.075 -13.135 ;
        RECT 94.250 -13.400 95.150 -13.385 ;
        RECT 96.245 -13.575 96.495 -12.975 ;
        RECT 93.590 -14.205 94.285 -13.575 ;
        RECT 96.165 -14.205 96.495 -13.575 ;
        RECT 36.150 -25.650 66.300 -25.250 ;
        RECT 26.300 -34.550 26.700 -32.750 ;
        RECT 30.050 -34.550 30.450 -32.750 ;
        RECT 31.850 -35.300 32.250 -32.750 ;
        RECT 33.950 -35.300 34.350 -32.700 ;
        RECT 34.650 -35.300 35.050 -32.750 ;
        RECT 31.850 -35.700 35.050 -35.300 ;
        RECT 35.550 -37.250 35.950 -32.750 ;
        RECT 36.450 -34.550 36.850 -32.750 ;
        RECT 37.350 -34.550 37.750 -32.750 ;
        RECT 39.450 -33.250 39.850 -32.750 ;
        RECT 40.150 -34.600 40.550 -32.800 ;
        RECT 41.050 -34.100 41.450 -32.800 ;
        RECT 43.000 -34.100 43.500 -26.450 ;
        RECT 47.315 -29.355 47.485 -28.595 ;
        RECT 47.315 -29.525 48.030 -29.355 ;
        RECT 48.200 -29.500 48.455 -28.595 ;
        RECT 47.225 -30.075 47.580 -29.705 ;
        RECT 47.860 -29.735 48.030 -29.525 ;
        RECT 47.860 -30.065 48.115 -29.735 ;
        RECT 47.860 -30.255 48.030 -30.065 ;
        RECT 48.285 -30.230 48.455 -29.500 ;
        RECT 47.315 -30.425 48.030 -30.255 ;
        RECT 47.315 -30.805 47.485 -30.425 ;
        RECT 48.200 -30.805 48.455 -30.230 ;
        RECT 55.455 -32.095 55.785 -31.295 ;
        RECT 56.295 -32.075 56.625 -31.295 ;
        RECT 59.665 -31.795 59.835 -31.295 ;
        RECT 59.665 -31.965 60.330 -31.795 ;
        RECT 56.295 -32.095 57.060 -32.075 ;
        RECT 55.455 -32.150 57.060 -32.095 ;
        RECT 59.580 -32.150 59.930 -32.135 ;
        RECT 55.455 -32.265 59.930 -32.150 ;
        RECT 54.995 -32.685 56.625 -32.435 ;
        RECT 56.795 -32.550 59.930 -32.265 ;
        RECT 56.795 -32.855 57.060 -32.550 ;
        RECT 59.580 -32.785 59.930 -32.550 ;
        RECT 55.455 -33.035 57.060 -32.855 ;
        RECT 60.100 -32.955 60.330 -31.965 ;
        RECT 55.455 -33.505 55.785 -33.035 ;
        RECT 56.295 -33.505 56.625 -33.035 ;
        RECT 58.100 -33.450 58.650 -33.000 ;
        RECT 59.665 -33.125 60.330 -32.955 ;
        RECT 59.665 -33.415 59.835 -33.125 ;
        RECT 60.505 -33.415 60.690 -31.295 ;
        RECT 61.365 -31.720 61.615 -31.295 ;
        RECT 61.825 -31.570 62.930 -31.400 ;
        RECT 61.310 -31.850 61.615 -31.720 ;
        RECT 60.860 -33.045 61.140 -32.095 ;
        RECT 61.310 -32.955 61.480 -31.850 ;
        RECT 61.650 -32.635 61.890 -32.040 ;
        RECT 62.060 -32.105 62.590 -31.740 ;
        RECT 62.060 -32.805 62.230 -32.105 ;
        RECT 62.760 -32.185 62.930 -31.570 ;
        RECT 63.440 -31.625 63.690 -31.295 ;
        RECT 63.915 -31.595 64.800 -31.425 ;
        RECT 62.760 -32.275 63.270 -32.185 ;
        RECT 61.310 -33.085 61.535 -32.955 ;
        RECT 61.705 -33.025 62.230 -32.805 ;
        RECT 62.400 -32.445 63.270 -32.275 ;
        RECT 61.365 -33.225 61.535 -33.085 ;
        RECT 62.400 -33.225 62.570 -32.445 ;
        RECT 63.100 -32.515 63.270 -32.445 ;
        RECT 62.780 -32.695 62.980 -32.665 ;
        RECT 63.440 -32.695 63.610 -31.625 ;
        RECT 63.780 -32.515 63.970 -31.795 ;
        RECT 62.780 -32.995 63.610 -32.695 ;
        RECT 64.140 -32.725 64.460 -31.765 ;
        RECT 61.365 -33.395 61.700 -33.225 ;
        RECT 61.895 -33.395 62.570 -33.225 ;
        RECT 63.440 -33.225 63.610 -32.995 ;
        RECT 63.995 -33.055 64.460 -32.725 ;
        RECT 64.630 -32.435 64.800 -31.595 ;
        RECT 65.525 -31.855 65.865 -31.295 ;
        RECT 64.970 -32.230 65.865 -31.855 ;
        RECT 65.675 -32.435 65.865 -32.230 ;
        RECT 66.375 -32.185 66.705 -31.340 ;
        RECT 66.375 -32.265 66.765 -32.185 ;
        RECT 66.550 -32.315 66.765 -32.265 ;
        RECT 64.630 -32.765 65.505 -32.435 ;
        RECT 65.675 -32.765 66.425 -32.435 ;
        RECT 64.630 -33.225 64.800 -32.765 ;
        RECT 65.675 -32.935 65.875 -32.765 ;
        RECT 66.595 -32.895 66.765 -32.315 ;
        RECT 66.540 -32.935 66.765 -32.895 ;
        RECT 63.440 -33.395 63.845 -33.225 ;
        RECT 64.015 -33.395 64.800 -33.225 ;
        RECT 41.050 -34.600 43.500 -34.100 ;
        RECT 58.275 -34.325 58.525 -33.450 ;
        RECT 65.545 -33.460 65.875 -32.935 ;
        RECT 66.385 -33.020 66.765 -32.935 ;
        RECT 66.385 -33.455 66.715 -33.020 ;
        RECT 27.450 -37.750 39.300 -37.250 ;
        RECT 27.450 -38.250 27.950 -37.750 ;
        RECT 25.050 -38.750 27.950 -38.250 ;
        RECT 25.050 -40.250 25.450 -38.750 ;
        RECT 18.595 -42.335 19.145 -42.165 ;
        RECT 18.975 -42.710 19.145 -42.335 ;
        RECT 19.325 -42.430 19.695 -42.075 ;
        RECT 19.875 -42.335 20.805 -42.165 ;
        RECT 19.875 -42.710 20.045 -42.335 ;
        RECT 18.975 -42.880 20.045 -42.710 ;
        RECT 19.335 -42.965 19.665 -42.880 ;
        RECT 18.595 -43.135 19.170 -43.050 ;
        RECT 19.900 -43.135 20.805 -43.050 ;
        RECT 18.595 -43.305 20.805 -43.135 ;
        RECT 19.450 -44.650 19.650 -43.305 ;
        RECT 25.750 -43.800 26.150 -39.800 ;
        RECT 26.150 -44.250 26.450 -44.200 ;
        RECT 21.850 -44.650 26.450 -44.250 ;
        RECT 19.450 -45.050 22.250 -44.650 ;
        RECT 26.150 -44.700 26.450 -44.650 ;
        RECT 19.450 -45.395 19.650 -45.050 ;
        RECT 19.415 -45.725 19.665 -45.395 ;
        RECT 26.650 -45.400 27.050 -39.800 ;
        RECT 27.550 -43.800 27.950 -38.750 ;
        RECT 27.250 -44.700 27.550 -44.200 ;
        RECT 30.550 -45.400 30.950 -39.950 ;
        RECT 31.450 -41.950 31.850 -37.750 ;
        RECT 32.350 -41.950 32.750 -39.950 ;
        RECT 34.400 -41.950 34.800 -39.950 ;
        RECT 35.300 -41.950 35.700 -37.750 ;
        RECT 38.900 -38.250 39.300 -37.750 ;
        RECT 38.900 -38.750 40.000 -38.250 ;
        RECT 31.150 -42.850 32.150 -42.350 ;
        RECT 35.100 -42.850 35.950 -42.350 ;
        RECT 26.650 -45.800 30.950 -45.400 ;
        RECT 18.595 -45.895 19.225 -45.815 ;
        RECT 19.825 -45.895 20.805 -45.815 ;
        RECT 18.595 -46.145 20.805 -45.895 ;
        RECT 31.450 -46.200 31.850 -42.850 ;
        RECT 36.200 -45.050 36.600 -39.950 ;
        RECT 38.900 -40.400 39.300 -38.750 ;
        RECT 39.600 -43.850 40.000 -38.750 ;
        RECT 40.000 -44.750 40.300 -44.250 ;
        RECT 40.500 -45.050 40.900 -39.850 ;
        RECT 41.400 -43.850 41.800 -39.850 ;
        RECT 41.100 -44.750 41.400 -44.250 ;
        RECT 43.000 -45.050 43.500 -34.600 ;
        RECT 57.500 -34.575 58.525 -34.325 ;
        RECT 52.785 -36.305 53.115 -35.495 ;
        RECT 52.785 -36.475 53.500 -36.305 ;
        RECT 52.780 -36.650 53.160 -36.645 ;
        RECT 51.200 -36.850 53.160 -36.650 ;
        RECT 51.200 -39.000 51.500 -36.850 ;
        RECT 52.780 -36.885 53.160 -36.850 ;
        RECT 53.330 -36.715 53.500 -36.475 ;
        RECT 53.705 -36.345 53.875 -35.495 ;
        RECT 54.545 -36.345 54.715 -35.495 ;
        RECT 57.500 -35.850 57.750 -34.575 ;
        RECT 53.705 -36.515 54.715 -36.345 ;
        RECT 54.220 -36.650 54.715 -36.515 ;
        RECT 55.450 -36.100 57.750 -35.850 ;
        RECT 58.265 -35.995 58.435 -35.495 ;
        RECT 55.450 -36.650 55.725 -36.100 ;
        RECT 58.265 -36.165 58.930 -35.995 ;
        RECT 53.330 -36.885 53.830 -36.715 ;
        RECT 53.330 -37.055 53.500 -36.885 ;
        RECT 54.220 -36.900 55.725 -36.650 ;
        RECT 54.220 -37.055 54.715 -36.900 ;
        RECT 58.180 -36.985 58.530 -36.335 ;
        RECT 52.865 -37.225 53.500 -37.055 ;
        RECT 53.705 -37.225 54.715 -37.055 ;
        RECT 58.700 -37.155 58.930 -36.165 ;
        RECT 52.865 -37.705 53.035 -37.225 ;
        RECT 53.705 -37.705 53.875 -37.225 ;
        RECT 54.545 -37.705 54.715 -37.225 ;
        RECT 58.265 -37.325 58.930 -37.155 ;
        RECT 58.265 -37.615 58.435 -37.325 ;
        RECT 59.105 -37.615 59.290 -35.495 ;
        RECT 59.965 -35.920 60.215 -35.495 ;
        RECT 60.425 -35.770 61.530 -35.600 ;
        RECT 59.910 -36.050 60.215 -35.920 ;
        RECT 59.460 -37.245 59.740 -36.295 ;
        RECT 59.910 -37.155 60.080 -36.050 ;
        RECT 60.250 -36.835 60.490 -36.240 ;
        RECT 60.660 -36.305 61.190 -35.940 ;
        RECT 60.660 -37.005 60.830 -36.305 ;
        RECT 61.360 -36.385 61.530 -35.770 ;
        RECT 62.040 -35.825 62.290 -35.495 ;
        RECT 62.515 -35.795 63.400 -35.625 ;
        RECT 61.360 -36.475 61.870 -36.385 ;
        RECT 59.910 -37.285 60.135 -37.155 ;
        RECT 60.305 -37.225 60.830 -37.005 ;
        RECT 61.000 -36.645 61.870 -36.475 ;
        RECT 59.965 -37.425 60.135 -37.285 ;
        RECT 61.000 -37.425 61.170 -36.645 ;
        RECT 61.700 -36.715 61.870 -36.645 ;
        RECT 61.380 -36.895 61.580 -36.865 ;
        RECT 62.040 -36.895 62.210 -35.825 ;
        RECT 62.380 -36.715 62.570 -35.995 ;
        RECT 61.380 -37.195 62.210 -36.895 ;
        RECT 62.740 -36.925 63.060 -35.965 ;
        RECT 59.965 -37.595 60.300 -37.425 ;
        RECT 60.495 -37.595 61.170 -37.425 ;
        RECT 62.040 -37.425 62.210 -37.195 ;
        RECT 62.595 -37.255 63.060 -36.925 ;
        RECT 63.230 -36.635 63.400 -35.795 ;
        RECT 64.130 -36.055 64.470 -35.495 ;
        RECT 63.570 -36.430 64.470 -36.055 ;
        RECT 64.280 -36.635 64.470 -36.430 ;
        RECT 64.980 -36.385 65.310 -35.540 ;
        RECT 65.995 -36.245 66.325 -35.515 ;
        RECT 64.980 -36.465 65.390 -36.385 ;
        RECT 65.155 -36.515 65.390 -36.465 ;
        RECT 63.230 -36.965 64.110 -36.635 ;
        RECT 64.280 -36.965 65.030 -36.635 ;
        RECT 63.230 -37.425 63.400 -36.965 ;
        RECT 64.280 -37.135 64.480 -36.965 ;
        RECT 65.200 -37.095 65.390 -36.515 ;
        RECT 65.145 -37.135 65.390 -37.095 ;
        RECT 62.040 -37.595 62.445 -37.425 ;
        RECT 62.615 -37.595 63.400 -37.425 ;
        RECT 64.150 -37.660 64.480 -37.135 ;
        RECT 64.990 -37.220 65.390 -37.135 ;
        RECT 66.055 -36.635 66.325 -36.245 ;
        RECT 66.900 -36.465 67.235 -35.495 ;
        RECT 78.315 -35.885 78.485 -35.125 ;
        RECT 66.055 -36.965 66.850 -36.635 ;
        RECT 67.020 -36.650 67.235 -36.465 ;
        RECT 74.200 -36.200 75.150 -36.000 ;
        RECT 78.315 -36.055 79.030 -35.885 ;
        RECT 79.200 -36.030 79.455 -35.125 ;
        RECT 81.755 -35.625 81.925 -35.125 ;
        RECT 81.755 -35.795 82.420 -35.625 ;
        RECT 74.200 -36.230 77.450 -36.200 ;
        RECT 74.200 -36.580 78.600 -36.230 ;
        RECT 78.860 -36.265 79.030 -36.055 ;
        RECT 74.200 -36.600 77.450 -36.580 ;
        RECT 67.020 -36.850 69.200 -36.650 ;
        RECT 64.990 -37.655 65.320 -37.220 ;
        RECT 66.055 -37.345 66.255 -36.965 ;
        RECT 67.020 -37.075 67.235 -36.850 ;
        RECT 67.850 -37.000 69.200 -36.850 ;
        RECT 74.200 -36.900 75.150 -36.600 ;
        RECT 78.225 -36.605 78.580 -36.580 ;
        RECT 78.860 -36.595 79.115 -36.265 ;
        RECT 79.285 -36.280 79.455 -36.030 ;
        RECT 81.670 -36.280 82.020 -35.965 ;
        RECT 79.285 -36.480 82.020 -36.280 ;
        RECT 78.860 -36.785 79.030 -36.595 ;
        RECT 79.285 -36.760 79.455 -36.480 ;
        RECT 81.670 -36.615 82.020 -36.480 ;
        RECT 65.995 -37.615 66.255 -37.345 ;
        RECT 66.980 -37.695 67.235 -37.075 ;
        RECT 68.000 -37.600 68.500 -37.200 ;
        RECT 68.800 -39.000 69.200 -37.000 ;
        RECT 78.315 -36.955 79.030 -36.785 ;
        RECT 78.315 -37.335 78.485 -36.955 ;
        RECT 79.200 -37.335 79.455 -36.760 ;
        RECT 82.190 -36.785 82.420 -35.795 ;
        RECT 81.755 -36.955 82.420 -36.785 ;
        RECT 81.755 -37.245 81.925 -36.955 ;
        RECT 82.595 -37.245 82.820 -35.125 ;
        RECT 83.535 -35.625 83.705 -35.125 ;
        RECT 83.940 -35.340 84.770 -35.170 ;
        RECT 83.010 -35.795 83.705 -35.625 ;
        RECT 83.010 -36.765 83.180 -35.795 ;
        RECT 83.350 -36.585 83.760 -35.965 ;
        RECT 83.930 -36.015 84.430 -35.635 ;
        RECT 83.010 -36.955 83.705 -36.765 ;
        RECT 83.930 -36.885 84.150 -36.015 ;
        RECT 84.600 -36.185 84.770 -35.340 ;
        RECT 85.570 -35.505 85.740 -35.215 ;
        RECT 86.710 -35.425 87.340 -35.175 ;
        RECT 87.170 -35.505 87.340 -35.425 ;
        RECT 88.140 -35.505 88.380 -35.215 ;
        RECT 84.940 -35.755 86.310 -35.505 ;
        RECT 84.940 -36.015 85.190 -35.755 ;
        RECT 85.700 -36.185 85.950 -36.025 ;
        RECT 84.600 -36.355 85.950 -36.185 ;
        RECT 84.600 -36.395 85.020 -36.355 ;
        RECT 84.330 -36.945 84.680 -36.575 ;
        RECT 83.535 -37.285 83.705 -36.955 ;
        RECT 84.850 -37.125 85.020 -36.395 ;
        RECT 86.120 -36.525 86.310 -35.755 ;
        RECT 85.190 -36.855 85.600 -36.525 ;
        RECT 84.005 -37.325 85.020 -37.125 ;
        RECT 85.890 -36.865 86.310 -36.525 ;
        RECT 86.480 -35.935 87.000 -35.625 ;
        RECT 87.170 -35.675 88.380 -35.505 ;
        RECT 86.480 -36.695 86.650 -35.935 ;
        RECT 86.820 -36.525 87.000 -36.115 ;
        RECT 87.170 -36.185 87.340 -35.675 ;
        RECT 89.110 -35.825 89.280 -35.215 ;
        RECT 89.550 -35.675 89.880 -35.165 ;
        RECT 89.110 -35.845 89.430 -35.825 ;
        RECT 87.510 -36.015 89.430 -35.845 ;
        RECT 87.170 -36.355 89.070 -36.185 ;
        RECT 87.400 -36.695 87.730 -36.575 ;
        RECT 86.480 -36.865 87.730 -36.695 ;
        RECT 85.890 -37.295 86.140 -36.865 ;
        RECT 87.900 -37.115 88.070 -36.355 ;
        RECT 88.740 -36.415 89.070 -36.355 ;
        RECT 88.260 -36.585 88.590 -36.525 ;
        RECT 88.260 -36.855 88.920 -36.585 ;
        RECT 89.240 -36.910 89.430 -36.015 ;
        RECT 87.220 -37.285 88.070 -37.115 ;
        RECT 89.110 -37.240 89.430 -36.910 ;
        RECT 89.630 -36.265 89.880 -35.675 ;
        RECT 90.525 -35.935 90.780 -35.265 ;
        RECT 90.600 -36.230 90.780 -35.935 ;
        RECT 93.225 -35.885 93.395 -35.125 ;
        RECT 93.225 -36.055 93.940 -35.885 ;
        RECT 94.110 -36.030 94.365 -35.125 ;
        RECT 90.600 -36.235 93.150 -36.230 ;
        RECT 89.630 -36.595 90.430 -36.265 ;
        RECT 89.630 -37.245 89.880 -36.595 ;
        RECT 90.600 -36.605 93.490 -36.235 ;
        RECT 93.770 -36.265 93.940 -36.055 ;
        RECT 93.770 -36.595 94.025 -36.265 ;
        RECT 90.600 -36.630 93.150 -36.605 ;
        RECT 90.600 -36.795 90.780 -36.630 ;
        RECT 93.770 -36.785 93.940 -36.595 ;
        RECT 94.195 -36.760 94.365 -36.030 ;
        RECT 90.525 -37.325 90.780 -36.795 ;
        RECT 93.225 -36.955 93.940 -36.785 ;
        RECT 93.225 -37.335 93.395 -36.955 ;
        RECT 94.110 -37.335 94.365 -36.760 ;
        RECT 51.200 -39.400 69.200 -39.000 ;
        RECT 78.815 -41.315 79.145 -40.335 ;
        RECT 78.895 -41.530 79.145 -41.315 ;
        RECT 86.385 -41.485 86.765 -40.805 ;
        RECT 87.695 -41.315 88.025 -40.805 ;
        RECT 88.535 -41.315 88.935 -40.805 ;
        RECT 87.695 -41.485 88.935 -41.315 ;
        RECT 78.895 -41.700 79.150 -41.530 ;
        RECT 78.895 -41.915 79.145 -41.700 ;
        RECT 78.815 -42.545 79.145 -41.915 ;
        RECT 86.385 -42.445 86.555 -41.485 ;
        RECT 86.725 -41.825 88.030 -41.655 ;
        RECT 89.115 -41.735 89.435 -40.805 ;
        RECT 91.055 -41.565 91.225 -40.805 ;
        RECT 91.055 -41.735 91.770 -41.565 ;
        RECT 91.940 -41.710 92.195 -40.805 ;
        RECT 86.725 -42.275 86.970 -41.825 ;
        RECT 87.140 -42.195 87.690 -41.995 ;
        RECT 87.860 -42.025 88.030 -41.825 ;
        RECT 88.805 -41.880 89.435 -41.735 ;
        RECT 88.805 -41.930 90.650 -41.880 ;
        RECT 90.965 -41.930 91.320 -41.915 ;
        RECT 87.860 -42.195 88.235 -42.025 ;
        RECT 88.405 -42.445 88.635 -41.945 ;
        RECT 86.385 -42.615 88.635 -42.445 ;
        RECT 88.805 -42.130 91.320 -41.930 ;
        RECT 86.935 -42.935 87.105 -42.615 ;
        RECT 88.805 -42.785 88.975 -42.130 ;
        RECT 90.965 -42.285 91.320 -42.130 ;
        RECT 91.600 -41.945 91.770 -41.735 ;
        RECT 91.600 -42.275 91.855 -41.945 ;
        RECT 91.600 -42.465 91.770 -42.275 ;
        RECT 92.025 -42.440 92.195 -41.710 ;
        RECT 88.020 -42.955 88.975 -42.785 ;
        RECT 91.055 -42.635 91.770 -42.465 ;
        RECT 55.455 -43.795 55.785 -42.995 ;
        RECT 56.295 -43.775 56.625 -42.995 ;
        RECT 59.665 -43.495 59.835 -42.995 ;
        RECT 59.665 -43.665 60.330 -43.495 ;
        RECT 56.295 -43.795 57.060 -43.775 ;
        RECT 55.455 -43.850 57.060 -43.795 ;
        RECT 59.580 -43.850 59.930 -43.835 ;
        RECT 55.455 -43.965 59.930 -43.850 ;
        RECT 54.995 -44.385 56.625 -44.135 ;
        RECT 56.795 -44.250 59.930 -43.965 ;
        RECT 56.795 -44.555 57.060 -44.250 ;
        RECT 59.580 -44.485 59.930 -44.250 ;
        RECT 36.200 -45.550 43.500 -45.050 ;
        RECT 55.455 -44.735 57.060 -44.555 ;
        RECT 60.100 -44.655 60.330 -43.665 ;
        RECT 55.455 -45.205 55.785 -44.735 ;
        RECT 56.295 -45.205 56.625 -44.735 ;
        RECT 58.100 -45.150 58.650 -44.700 ;
        RECT 59.665 -44.825 60.330 -44.655 ;
        RECT 59.665 -45.115 59.835 -44.825 ;
        RECT 60.505 -45.115 60.690 -42.995 ;
        RECT 61.365 -43.420 61.615 -42.995 ;
        RECT 61.825 -43.270 62.930 -43.100 ;
        RECT 61.310 -43.550 61.615 -43.420 ;
        RECT 60.860 -44.745 61.140 -43.795 ;
        RECT 61.310 -44.655 61.480 -43.550 ;
        RECT 61.650 -44.335 61.890 -43.740 ;
        RECT 62.060 -43.805 62.590 -43.440 ;
        RECT 62.060 -44.505 62.230 -43.805 ;
        RECT 62.760 -43.885 62.930 -43.270 ;
        RECT 63.440 -43.325 63.690 -42.995 ;
        RECT 63.915 -43.295 64.800 -43.125 ;
        RECT 62.760 -43.975 63.270 -43.885 ;
        RECT 61.310 -44.785 61.535 -44.655 ;
        RECT 61.705 -44.725 62.230 -44.505 ;
        RECT 62.400 -44.145 63.270 -43.975 ;
        RECT 61.365 -44.925 61.535 -44.785 ;
        RECT 62.400 -44.925 62.570 -44.145 ;
        RECT 63.100 -44.215 63.270 -44.145 ;
        RECT 62.780 -44.395 62.980 -44.365 ;
        RECT 63.440 -44.395 63.610 -43.325 ;
        RECT 63.780 -44.215 63.970 -43.495 ;
        RECT 62.780 -44.695 63.610 -44.395 ;
        RECT 64.140 -44.425 64.460 -43.465 ;
        RECT 61.365 -45.095 61.700 -44.925 ;
        RECT 61.895 -45.095 62.570 -44.925 ;
        RECT 63.440 -44.925 63.610 -44.695 ;
        RECT 63.995 -44.755 64.460 -44.425 ;
        RECT 64.630 -44.135 64.800 -43.295 ;
        RECT 65.525 -43.555 65.865 -42.995 ;
        RECT 91.055 -43.015 91.225 -42.635 ;
        RECT 91.940 -43.015 92.195 -42.440 ;
        RECT 64.970 -43.930 65.865 -43.555 ;
        RECT 65.675 -44.135 65.865 -43.930 ;
        RECT 66.375 -43.885 66.705 -43.040 ;
        RECT 66.375 -43.965 66.765 -43.885 ;
        RECT 66.550 -44.015 66.765 -43.965 ;
        RECT 64.630 -44.465 65.505 -44.135 ;
        RECT 65.675 -44.465 66.425 -44.135 ;
        RECT 64.630 -44.925 64.800 -44.465 ;
        RECT 65.675 -44.635 65.875 -44.465 ;
        RECT 66.595 -44.595 66.765 -44.015 ;
        RECT 66.540 -44.635 66.765 -44.595 ;
        RECT 63.440 -45.095 63.845 -44.925 ;
        RECT 64.015 -45.095 64.800 -44.925 ;
        RECT 58.275 -46.025 58.525 -45.150 ;
        RECT 65.545 -45.160 65.875 -44.635 ;
        RECT 66.385 -44.720 66.765 -44.635 ;
        RECT 66.385 -45.155 66.715 -44.720 ;
        RECT 21.850 -46.700 41.800 -46.200 ;
        RECT 57.500 -46.275 58.525 -46.025 ;
        RECT 79.675 -46.125 80.005 -45.495 ;
        RECT 82.080 -46.035 82.335 -45.505 ;
        RECT 21.850 -47.300 22.350 -46.700 ;
        RECT 19.700 -47.800 22.350 -47.300 ;
        RECT 52.785 -48.005 53.115 -47.195 ;
        RECT 52.785 -48.175 53.500 -48.005 ;
        RECT 52.780 -48.350 53.160 -48.345 ;
        RECT 51.200 -48.550 53.160 -48.350 ;
        RECT 27.930 -49.520 30.090 -49.170 ;
        RECT 51.200 -50.700 51.500 -48.550 ;
        RECT 52.780 -48.585 53.160 -48.550 ;
        RECT 53.330 -48.415 53.500 -48.175 ;
        RECT 53.705 -48.045 53.875 -47.195 ;
        RECT 54.545 -48.045 54.715 -47.195 ;
        RECT 57.500 -47.550 57.750 -46.275 ;
        RECT 79.675 -46.725 79.925 -46.125 ;
        RECT 80.095 -46.320 80.425 -46.315 ;
        RECT 82.080 -46.320 82.260 -46.035 ;
        RECT 82.980 -46.235 83.230 -45.585 ;
        RECT 80.095 -46.560 82.260 -46.320 ;
        RECT 80.095 -46.565 80.425 -46.560 ;
        RECT 53.705 -48.215 54.715 -48.045 ;
        RECT 54.220 -48.350 54.715 -48.215 ;
        RECT 55.450 -47.800 57.750 -47.550 ;
        RECT 58.265 -47.695 58.435 -47.195 ;
        RECT 55.450 -48.350 55.725 -47.800 ;
        RECT 58.265 -47.865 58.930 -47.695 ;
        RECT 53.330 -48.585 53.830 -48.415 ;
        RECT 53.330 -48.755 53.500 -48.585 ;
        RECT 54.220 -48.600 55.725 -48.350 ;
        RECT 54.220 -48.755 54.715 -48.600 ;
        RECT 58.180 -48.685 58.530 -48.035 ;
        RECT 52.865 -48.925 53.500 -48.755 ;
        RECT 53.705 -48.925 54.715 -48.755 ;
        RECT 58.700 -48.855 58.930 -47.865 ;
        RECT 52.865 -49.405 53.035 -48.925 ;
        RECT 53.705 -49.405 53.875 -48.925 ;
        RECT 54.545 -49.405 54.715 -48.925 ;
        RECT 58.265 -49.025 58.930 -48.855 ;
        RECT 58.265 -49.315 58.435 -49.025 ;
        RECT 59.105 -49.315 59.290 -47.195 ;
        RECT 59.965 -47.620 60.215 -47.195 ;
        RECT 60.425 -47.470 61.530 -47.300 ;
        RECT 59.910 -47.750 60.215 -47.620 ;
        RECT 59.460 -48.945 59.740 -47.995 ;
        RECT 59.910 -48.855 60.080 -47.750 ;
        RECT 60.250 -48.535 60.490 -47.940 ;
        RECT 60.660 -48.005 61.190 -47.640 ;
        RECT 60.660 -48.705 60.830 -48.005 ;
        RECT 61.360 -48.085 61.530 -47.470 ;
        RECT 62.040 -47.525 62.290 -47.195 ;
        RECT 62.515 -47.495 63.400 -47.325 ;
        RECT 61.360 -48.175 61.870 -48.085 ;
        RECT 59.910 -48.985 60.135 -48.855 ;
        RECT 60.305 -48.925 60.830 -48.705 ;
        RECT 61.000 -48.345 61.870 -48.175 ;
        RECT 59.965 -49.125 60.135 -48.985 ;
        RECT 61.000 -49.125 61.170 -48.345 ;
        RECT 61.700 -48.415 61.870 -48.345 ;
        RECT 61.380 -48.595 61.580 -48.565 ;
        RECT 62.040 -48.595 62.210 -47.525 ;
        RECT 62.380 -48.415 62.570 -47.695 ;
        RECT 61.380 -48.895 62.210 -48.595 ;
        RECT 62.740 -48.625 63.060 -47.665 ;
        RECT 59.965 -49.295 60.300 -49.125 ;
        RECT 60.495 -49.295 61.170 -49.125 ;
        RECT 62.040 -49.125 62.210 -48.895 ;
        RECT 62.595 -48.955 63.060 -48.625 ;
        RECT 63.230 -48.335 63.400 -47.495 ;
        RECT 64.130 -47.755 64.470 -47.195 ;
        RECT 63.570 -48.130 64.470 -47.755 ;
        RECT 64.280 -48.335 64.470 -48.130 ;
        RECT 64.980 -48.085 65.310 -47.240 ;
        RECT 65.995 -47.945 66.325 -47.215 ;
        RECT 64.980 -48.165 65.390 -48.085 ;
        RECT 65.155 -48.215 65.390 -48.165 ;
        RECT 63.230 -48.665 64.110 -48.335 ;
        RECT 64.280 -48.665 65.030 -48.335 ;
        RECT 63.230 -49.125 63.400 -48.665 ;
        RECT 64.280 -48.835 64.480 -48.665 ;
        RECT 65.200 -48.795 65.390 -48.215 ;
        RECT 65.145 -48.835 65.390 -48.795 ;
        RECT 62.040 -49.295 62.445 -49.125 ;
        RECT 62.615 -49.295 63.400 -49.125 ;
        RECT 64.150 -49.360 64.480 -48.835 ;
        RECT 64.990 -48.920 65.390 -48.835 ;
        RECT 66.055 -48.335 66.325 -47.945 ;
        RECT 66.900 -48.165 67.235 -47.195 ;
        RECT 79.675 -47.705 80.005 -46.725 ;
        RECT 82.080 -46.895 82.260 -46.560 ;
        RECT 82.430 -46.565 83.230 -46.235 ;
        RECT 82.080 -47.565 82.335 -46.895 ;
        RECT 82.980 -47.155 83.230 -46.565 ;
        RECT 83.430 -45.920 83.750 -45.590 ;
        RECT 84.790 -45.715 85.640 -45.545 ;
        RECT 83.430 -46.815 83.620 -45.920 ;
        RECT 83.940 -46.245 84.600 -45.975 ;
        RECT 84.270 -46.305 84.600 -46.245 ;
        RECT 83.790 -46.475 84.120 -46.415 ;
        RECT 84.790 -46.475 84.960 -45.715 ;
        RECT 86.720 -45.965 86.970 -45.535 ;
        RECT 85.130 -46.135 86.380 -45.965 ;
        RECT 85.130 -46.255 85.460 -46.135 ;
        RECT 83.790 -46.645 85.690 -46.475 ;
        RECT 83.430 -46.985 85.350 -46.815 ;
        RECT 83.430 -47.005 83.750 -46.985 ;
        RECT 82.980 -47.665 83.310 -47.155 ;
        RECT 83.580 -47.615 83.750 -47.005 ;
        RECT 85.520 -47.155 85.690 -46.645 ;
        RECT 85.860 -46.715 86.040 -46.305 ;
        RECT 86.210 -46.895 86.380 -46.135 ;
        RECT 84.480 -47.325 85.690 -47.155 ;
        RECT 85.860 -47.205 86.380 -46.895 ;
        RECT 86.550 -46.305 86.970 -45.965 ;
        RECT 87.840 -45.705 88.855 -45.505 ;
        RECT 87.260 -46.305 87.670 -45.975 ;
        RECT 86.550 -47.075 86.740 -46.305 ;
        RECT 87.840 -46.435 88.010 -45.705 ;
        RECT 89.155 -45.875 89.325 -45.545 ;
        RECT 88.180 -46.255 88.530 -45.885 ;
        RECT 87.840 -46.475 88.260 -46.435 ;
        RECT 86.910 -46.645 88.260 -46.475 ;
        RECT 86.910 -46.805 87.160 -46.645 ;
        RECT 87.670 -47.075 87.920 -46.815 ;
        RECT 86.550 -47.325 87.920 -47.075 ;
        RECT 84.480 -47.615 84.720 -47.325 ;
        RECT 85.520 -47.405 85.690 -47.325 ;
        RECT 85.520 -47.655 86.150 -47.405 ;
        RECT 87.120 -47.615 87.290 -47.325 ;
        RECT 88.090 -47.490 88.260 -46.645 ;
        RECT 88.710 -46.815 88.930 -45.945 ;
        RECT 89.155 -46.065 89.850 -45.875 ;
        RECT 88.430 -47.195 88.930 -46.815 ;
        RECT 89.100 -46.865 89.510 -46.245 ;
        RECT 89.680 -47.035 89.850 -46.065 ;
        RECT 89.155 -47.205 89.850 -47.035 ;
        RECT 88.090 -47.660 88.920 -47.490 ;
        RECT 89.155 -47.705 89.325 -47.205 ;
        RECT 90.040 -47.705 90.265 -45.585 ;
        RECT 90.935 -45.875 91.105 -45.585 ;
        RECT 90.440 -46.045 91.105 -45.875 ;
        RECT 90.440 -47.035 90.670 -46.045 ;
        RECT 93.735 -46.070 93.990 -45.495 ;
        RECT 94.705 -45.875 94.875 -45.495 ;
        RECT 94.160 -46.045 94.875 -45.875 ;
        RECT 90.840 -46.230 91.190 -46.215 ;
        RECT 90.840 -46.580 92.750 -46.230 ;
        RECT 90.840 -46.865 91.190 -46.580 ;
        RECT 93.735 -46.800 93.905 -46.070 ;
        RECT 94.160 -46.235 94.330 -46.045 ;
        RECT 95.400 -46.180 95.900 -46.150 ;
        RECT 95.250 -46.220 95.900 -46.180 ;
        RECT 94.075 -46.565 94.330 -46.235 ;
        RECT 94.160 -46.775 94.330 -46.565 ;
        RECT 94.610 -46.600 95.900 -46.220 ;
        RECT 95.250 -46.630 95.900 -46.600 ;
        RECT 95.400 -46.650 95.900 -46.630 ;
        RECT 90.440 -47.205 91.105 -47.035 ;
        RECT 90.935 -47.705 91.105 -47.205 ;
        RECT 93.735 -47.705 93.990 -46.800 ;
        RECT 94.160 -46.945 94.875 -46.775 ;
        RECT 94.705 -47.705 94.875 -46.945 ;
        RECT 66.055 -48.665 66.850 -48.335 ;
        RECT 67.020 -48.350 67.235 -48.165 ;
        RECT 67.020 -48.550 69.200 -48.350 ;
        RECT 64.990 -49.355 65.320 -48.920 ;
        RECT 66.055 -49.045 66.255 -48.665 ;
        RECT 67.020 -48.775 67.235 -48.550 ;
        RECT 67.850 -48.700 69.200 -48.550 ;
        RECT 65.995 -49.315 66.255 -49.045 ;
        RECT 66.980 -49.395 67.235 -48.775 ;
        RECT 68.000 -49.300 68.500 -48.900 ;
        RECT 68.800 -50.700 69.200 -48.700 ;
        RECT 51.200 -51.100 69.200 -50.700 ;
      LAYER met1 ;
        RECT -2.150 35.650 -1.750 36.150 ;
        RECT 12.800 35.650 13.200 36.150 ;
        RECT 27.850 35.650 28.250 36.150 ;
        RECT 42.800 35.650 43.200 36.150 ;
        RECT 57.850 35.650 58.250 36.150 ;
        RECT 72.800 35.650 73.200 36.150 ;
        RECT -10.100 35.150 -3.100 35.650 ;
        RECT -10.100 8.300 -9.600 35.150 ;
        RECT -3.600 32.050 -3.100 35.150 ;
        RECT -2.150 35.150 26.900 35.650 ;
        RECT -2.150 34.750 -1.750 35.150 ;
        RECT 5.200 32.050 5.700 35.150 ;
        RECT 12.800 34.750 13.200 35.150 ;
        RECT 7.350 34.100 7.750 34.450 ;
        RECT 18.250 34.100 18.650 34.450 ;
        RECT 7.350 33.600 18.650 34.100 ;
        RECT 7.350 33.250 7.750 33.600 ;
        RECT 10.050 32.050 10.550 33.600 ;
        RECT 18.250 33.250 18.650 33.600 ;
        RECT 26.400 32.050 26.900 35.150 ;
        RECT 27.850 35.150 56.900 35.650 ;
        RECT 27.850 34.750 28.250 35.150 ;
        RECT 35.200 32.050 35.700 35.150 ;
        RECT 42.800 34.750 43.200 35.150 ;
        RECT 37.350 34.100 37.750 34.450 ;
        RECT 48.250 34.100 48.650 34.450 ;
        RECT 37.350 33.600 48.650 34.100 ;
        RECT 37.350 33.250 37.750 33.600 ;
        RECT 40.050 32.050 40.550 33.600 ;
        RECT 48.250 33.250 48.650 33.600 ;
        RECT 56.400 32.050 56.900 35.150 ;
        RECT 57.850 35.150 85.900 35.650 ;
        RECT 57.850 34.750 58.250 35.150 ;
        RECT 65.200 32.050 65.700 35.150 ;
        RECT 72.800 34.750 73.200 35.150 ;
        RECT 67.350 34.100 67.750 34.450 ;
        RECT 78.250 34.100 78.650 34.450 ;
        RECT 67.350 33.600 78.650 34.100 ;
        RECT 67.350 33.250 67.750 33.600 ;
        RECT 70.050 32.050 70.550 33.600 ;
        RECT 78.250 33.250 78.650 33.600 ;
        RECT -5.000 31.400 -0.100 32.050 ;
        RECT 4.850 31.400 6.050 32.050 ;
        RECT 9.700 31.400 10.900 32.050 ;
        RECT 15.400 31.950 20.300 32.050 ;
        RECT 14.550 31.450 20.300 31.950 ;
        RECT 14.550 29.300 15.050 31.450 ;
        RECT 15.400 31.400 20.300 31.450 ;
        RECT 25.000 31.400 29.900 32.050 ;
        RECT 34.850 31.400 36.050 32.050 ;
        RECT 39.700 31.400 40.900 32.050 ;
        RECT 45.400 31.950 50.300 32.050 ;
        RECT 44.550 31.450 50.300 31.950 ;
        RECT -8.600 28.800 15.050 29.300 ;
        RECT 18.250 29.300 18.650 29.600 ;
        RECT 44.550 29.300 45.050 31.450 ;
        RECT 45.400 31.400 50.300 31.450 ;
        RECT 55.000 31.400 59.900 32.050 ;
        RECT 64.850 31.400 66.050 32.050 ;
        RECT 69.700 31.400 70.900 32.050 ;
        RECT 75.400 31.950 80.300 32.050 ;
        RECT 74.550 31.450 80.300 31.950 ;
        RECT 18.250 28.800 45.050 29.300 ;
        RECT 48.250 29.300 48.650 29.600 ;
        RECT 74.550 29.300 75.050 31.450 ;
        RECT 75.400 31.400 80.300 31.450 ;
        RECT 48.250 28.800 75.050 29.300 ;
        RECT 78.250 29.300 78.650 29.600 ;
        RECT 78.250 28.800 84.400 29.300 ;
        RECT -8.600 14.650 -8.100 28.800 ;
        RECT 18.250 28.400 18.650 28.800 ;
        RECT 48.250 28.400 48.650 28.800 ;
        RECT 78.250 28.400 78.650 28.800 ;
        RECT 14.825 22.450 16.930 22.830 ;
        RECT 24.970 20.900 27.075 21.280 ;
        RECT 17.300 17.400 17.750 17.500 ;
        RECT 14.350 17.100 17.750 17.400 ;
        RECT 14.350 14.650 14.850 17.100 ;
        RECT 17.300 17.050 17.750 17.100 ;
        RECT 27.150 14.650 27.550 15.050 ;
        RECT 57.150 14.650 57.550 15.050 ;
        RECT 83.900 14.650 84.400 28.800 ;
        RECT -8.600 14.150 27.550 14.650 ;
        RECT 27.150 13.850 27.550 14.150 ;
        RECT 30.750 14.150 57.550 14.650 ;
        RECT 25.500 12.000 30.400 12.050 ;
        RECT 30.750 12.000 31.250 14.150 ;
        RECT 57.150 13.850 57.550 14.150 ;
        RECT 60.750 14.150 84.400 14.650 ;
        RECT 25.500 11.500 31.250 12.000 ;
        RECT 25.500 11.400 30.400 11.500 ;
        RECT 34.900 11.400 36.100 12.050 ;
        RECT 39.750 11.400 40.950 12.050 ;
        RECT 45.900 11.400 50.800 12.050 ;
        RECT 55.500 12.000 60.400 12.050 ;
        RECT 60.750 12.000 61.250 14.150 ;
        RECT 55.500 11.500 61.250 12.000 ;
        RECT 55.500 11.400 60.400 11.500 ;
        RECT 64.900 11.400 66.100 12.050 ;
        RECT 69.750 11.400 70.950 12.050 ;
        RECT 75.900 11.400 80.800 12.050 ;
        RECT 27.150 9.850 27.550 10.200 ;
        RECT 35.250 9.850 35.750 11.400 ;
        RECT 38.050 9.850 38.450 10.200 ;
        RECT 27.150 9.350 38.450 9.850 ;
        RECT 27.150 9.000 27.550 9.350 ;
        RECT 38.050 9.000 38.450 9.350 ;
        RECT 32.600 8.300 33.000 8.700 ;
        RECT 40.100 8.300 40.600 11.400 ;
        RECT 47.550 8.300 47.950 8.700 ;
        RECT -16.950 7.800 47.950 8.300 ;
        RECT 48.900 8.300 49.400 11.400 ;
        RECT 57.150 9.850 57.550 10.200 ;
        RECT 65.250 9.850 65.750 11.400 ;
        RECT 68.050 9.850 68.450 10.200 ;
        RECT 57.150 9.350 68.450 9.850 ;
        RECT 57.150 9.000 57.550 9.350 ;
        RECT 68.050 9.000 68.450 9.350 ;
        RECT 62.600 8.300 63.000 8.700 ;
        RECT 70.100 8.300 70.600 11.400 ;
        RECT 77.550 8.300 77.950 8.700 ;
        RECT 48.900 7.800 77.950 8.300 ;
        RECT 78.900 8.300 79.400 11.400 ;
        RECT 85.400 8.300 85.900 35.150 ;
        RECT 78.900 7.800 85.900 8.300 ;
        RECT -16.950 -14.150 -16.500 7.800 ;
        RECT 32.600 7.300 33.000 7.800 ;
        RECT 47.550 7.300 47.950 7.800 ;
        RECT 62.600 7.300 63.000 7.800 ;
        RECT 77.550 7.300 77.950 7.800 ;
        RECT 21.700 -3.850 68.700 -3.450 ;
        RECT 21.700 -6.400 22.100 -3.850 ;
        RECT 26.000 -6.500 26.400 -3.850 ;
        RECT 28.900 -6.500 29.300 -3.850 ;
        RECT 31.800 -6.400 32.200 -3.850 ;
        RECT 36.100 -6.400 36.500 -3.850 ;
        RECT 40.400 -6.500 40.800 -3.850 ;
        RECT 43.300 -6.500 43.700 -3.850 ;
        RECT 46.200 -6.400 46.600 -3.850 ;
        RECT 50.500 -6.400 50.900 -3.850 ;
        RECT 54.800 -6.500 55.200 -3.850 ;
        RECT 57.700 -6.500 58.100 -3.850 ;
        RECT 60.600 -6.400 61.000 -3.850 ;
        RECT 23.800 -6.950 24.200 -6.750 ;
        RECT 31.000 -6.950 31.400 -6.750 ;
        RECT 23.800 -7.150 31.400 -6.950 ;
        RECT 38.200 -6.950 38.600 -6.750 ;
        RECT 45.400 -6.950 45.800 -6.750 ;
        RECT 38.200 -7.150 45.800 -6.950 ;
        RECT 52.600 -6.950 53.000 -6.750 ;
        RECT 59.800 -6.950 60.200 -6.750 ;
        RECT 52.600 -7.150 60.200 -6.950 ;
        RECT 19.000 -7.550 23.450 -7.150 ;
        RECT 23.800 -7.350 37.850 -7.150 ;
        RECT 23.800 -7.550 24.200 -7.350 ;
        RECT -11.220 -13.600 -10.930 -13.555 ;
        RECT -9.360 -13.600 -9.070 -13.555 ;
        RECT -6.580 -13.600 -6.290 -13.555 ;
        RECT -11.220 -13.740 -6.290 -13.600 ;
        RECT -11.220 -13.785 -10.930 -13.740 ;
        RECT -9.360 -13.785 -9.070 -13.740 ;
        RECT -6.580 -13.785 -6.290 -13.740 ;
        RECT 0.750 -13.780 3.050 -13.430 ;
        RECT -16.950 -14.600 -16.000 -14.150 ;
        RECT -12.750 -14.430 -9.600 -14.030 ;
        RECT -6.580 -14.280 -6.290 -14.235 ;
        RECT -8.825 -14.420 -6.290 -14.280 ;
        RECT -14.050 -19.380 -13.600 -19.330 ;
        RECT -14.450 -19.730 -13.600 -19.380 ;
        RECT -14.050 -19.780 -13.600 -19.730 ;
        RECT -12.750 -21.280 -12.400 -14.430 ;
        RECT -8.825 -14.575 -8.610 -14.420 ;
        RECT -6.580 -14.465 -6.290 -14.420 ;
        RECT -10.760 -14.620 -10.470 -14.575 ;
        RECT -8.900 -14.620 -8.610 -14.575 ;
        RECT -7.980 -14.580 -7.690 -14.575 ;
        RECT -10.760 -14.760 -8.610 -14.620 ;
        RECT -10.760 -14.805 -10.470 -14.760 ;
        RECT -8.900 -14.805 -8.610 -14.760 ;
        RECT -8.050 -14.620 -7.550 -14.580 ;
        RECT -4.720 -14.620 -4.430 -14.575 ;
        RECT -8.050 -14.760 -4.430 -14.620 ;
        RECT -8.050 -15.030 -7.550 -14.760 ;
        RECT -4.720 -14.805 -4.430 -14.760 ;
        RECT -1.300 -17.030 -0.950 -14.180 ;
        RECT -8.650 -17.380 -0.950 -17.030 ;
        RECT -8.650 -19.030 -8.300 -17.380 ;
        RECT -8.650 -19.380 -5.750 -19.030 ;
        RECT -6.700 -20.230 -6.350 -19.880 ;
        RECT -6.100 -19.930 -5.750 -19.380 ;
        RECT -1.450 -19.830 -1.150 -19.130 ;
        RECT -0.350 -19.830 0.300 -19.800 ;
        RECT -6.200 -20.180 -5.650 -19.930 ;
        RECT -1.450 -20.180 0.300 -19.830 ;
        RECT -1.450 -20.190 -1.150 -20.180 ;
        RECT -0.350 -20.200 0.300 -20.180 ;
        RECT -15.400 -21.580 -12.400 -21.280 ;
        RECT -8.650 -20.580 -6.350 -20.230 ;
        RECT -15.400 -23.730 -15.050 -21.580 ;
        RECT -8.650 -22.280 -8.300 -20.580 ;
        RECT 2.700 -22.080 3.050 -13.780 ;
        RECT -12.400 -22.630 -8.300 -22.280 ;
        RECT -1.650 -22.430 3.050 -22.080 ;
        RECT -12.400 -23.680 -12.050 -22.630 ;
        RECT -15.400 -24.080 -13.350 -23.730 ;
        RECT -12.400 -24.080 -10.950 -23.680 ;
        RECT -9.410 -23.970 -9.120 -23.925 ;
        RECT -6.150 -23.970 -5.650 -23.630 ;
        RECT -9.410 -24.110 -5.650 -23.970 ;
        RECT -9.410 -24.155 -9.120 -24.110 ;
        RECT -6.150 -24.130 -5.650 -24.110 ;
        RECT -5.230 -23.970 -4.940 -23.925 ;
        RECT -3.370 -23.970 -3.080 -23.925 ;
        RECT -5.230 -24.110 -3.080 -23.970 ;
        RECT -6.150 -24.155 -5.860 -24.130 ;
        RECT -5.230 -24.155 -4.940 -24.110 ;
        RECT -3.370 -24.155 -3.080 -24.110 ;
        RECT -7.550 -24.310 -7.260 -24.265 ;
        RECT -5.230 -24.310 -5.015 -24.155 ;
        RECT -7.550 -24.450 -5.015 -24.310 ;
        RECT -7.550 -24.495 -7.260 -24.450 ;
        RECT -4.250 -24.480 -3.850 -24.280 ;
        RECT -1.650 -24.480 -1.300 -22.430 ;
        RECT 19.000 -22.750 19.500 -7.550 ;
        RECT 23.050 -9.300 23.450 -7.550 ;
        RECT 23.050 -9.750 24.900 -9.300 ;
        RECT 27.350 -9.700 27.750 -7.350 ;
        RECT 31.000 -7.550 37.850 -7.350 ;
        RECT 38.200 -7.350 52.250 -7.150 ;
        RECT 38.200 -7.550 38.600 -7.350 ;
        RECT 31.000 -7.950 31.400 -7.550 ;
        RECT 28.100 -8.750 34.300 -8.350 ;
        RECT 30.250 -9.700 30.650 -8.750 ;
        RECT 37.450 -9.300 37.850 -7.550 ;
        RECT 33.150 -9.750 35.000 -9.300 ;
        RECT 37.450 -9.750 39.300 -9.300 ;
        RECT 41.750 -9.700 42.150 -7.350 ;
        RECT 45.400 -7.550 52.250 -7.350 ;
        RECT 52.600 -7.350 67.200 -7.150 ;
        RECT 52.600 -7.550 53.000 -7.350 ;
        RECT 45.400 -7.950 45.800 -7.550 ;
        RECT 42.500 -8.750 48.700 -8.350 ;
        RECT 44.650 -9.700 45.050 -8.750 ;
        RECT 51.850 -9.300 52.250 -7.550 ;
        RECT 47.550 -9.750 49.400 -9.300 ;
        RECT 51.850 -9.750 53.700 -9.300 ;
        RECT 56.150 -9.700 56.550 -7.350 ;
        RECT 59.800 -7.550 67.200 -7.350 ;
        RECT 59.800 -7.950 60.200 -7.550 ;
        RECT 56.900 -8.750 63.100 -8.350 ;
        RECT 59.050 -9.700 59.450 -8.750 ;
        RECT 61.950 -9.750 63.800 -9.300 ;
        RECT 33.150 -10.850 33.600 -9.750 ;
        RECT 20.500 -11.250 33.600 -10.850 ;
        RECT 33.900 -10.850 34.300 -10.450 ;
        RECT 47.550 -10.850 48.000 -9.750 ;
        RECT 33.900 -11.250 48.000 -10.850 ;
        RECT 48.300 -10.850 48.700 -10.450 ;
        RECT 61.950 -10.850 62.400 -9.750 ;
        RECT 48.300 -11.250 62.400 -10.850 ;
        RECT 62.700 -10.850 63.100 -10.450 ;
        RECT 62.700 -11.250 65.700 -10.850 ;
        RECT 20.500 -19.050 21.000 -11.250 ;
        RECT 33.900 -11.650 34.300 -11.250 ;
        RECT 48.300 -11.650 48.700 -11.250 ;
        RECT 62.700 -11.650 63.100 -11.250 ;
        RECT 37.550 -19.050 37.950 -18.650 ;
        RECT 51.950 -19.050 52.350 -18.650 ;
        RECT 65.200 -19.050 65.700 -11.250 ;
        RECT 20.500 -19.450 37.950 -19.050 ;
        RECT 37.550 -19.850 37.950 -19.450 ;
        RECT 38.250 -19.450 52.350 -19.050 ;
        RECT 38.250 -20.550 38.700 -19.450 ;
        RECT 51.950 -19.850 52.350 -19.450 ;
        RECT 52.650 -19.450 65.700 -19.050 ;
        RECT 52.650 -20.550 53.100 -19.450 ;
        RECT 36.850 -21.000 38.700 -20.550 ;
        RECT 41.200 -21.550 41.600 -20.600 ;
        RECT 37.550 -21.950 43.750 -21.550 ;
        RECT 40.450 -22.750 40.850 -22.350 ;
        RECT 19.000 -22.950 40.850 -22.750 ;
        RECT 44.100 -22.950 44.500 -20.600 ;
        RECT 46.950 -21.000 48.800 -20.550 ;
        RECT 51.250 -21.000 53.100 -20.550 ;
        RECT 48.400 -22.750 48.800 -21.000 ;
        RECT 55.600 -21.550 56.000 -20.600 ;
        RECT 51.950 -21.950 58.150 -21.550 ;
        RECT 54.850 -22.750 55.250 -22.350 ;
        RECT 47.650 -22.950 48.050 -22.750 ;
        RECT 19.000 -23.150 48.050 -22.950 ;
        RECT 48.400 -22.950 55.250 -22.750 ;
        RECT 58.500 -22.950 58.900 -20.600 ;
        RECT 61.350 -21.000 63.200 -20.550 ;
        RECT 62.800 -22.750 63.200 -21.000 ;
        RECT 66.700 -22.750 67.200 -7.550 ;
        RECT 62.050 -22.950 62.450 -22.750 ;
        RECT 48.400 -23.150 62.450 -22.950 ;
        RECT 62.800 -23.150 67.200 -22.750 ;
        RECT -4.250 -24.780 -1.300 -24.480 ;
        RECT -0.950 -24.530 0.700 -24.180 ;
        RECT -4.250 -24.830 -3.050 -24.780 ;
        RECT -2.450 -24.830 -1.300 -24.780 ;
        RECT -7.550 -24.990 -7.260 -24.945 ;
        RECT -4.770 -24.990 -4.480 -24.945 ;
        RECT -2.910 -24.990 -2.620 -24.945 ;
        RECT -7.550 -25.130 -2.620 -24.990 ;
        RECT -7.550 -25.175 -7.260 -25.130 ;
        RECT -4.770 -25.175 -4.480 -25.130 ;
        RECT -2.910 -25.175 -2.620 -25.130 ;
        RECT 0.350 -25.330 0.700 -24.530 ;
        RECT 2.350 -62.450 2.850 -24.100 ;
        RECT 34.200 -28.050 34.600 -23.150 ;
        RECT 40.450 -23.350 48.050 -23.150 ;
        RECT 40.450 -23.550 40.850 -23.350 ;
        RECT 47.650 -23.550 48.050 -23.350 ;
        RECT 54.850 -23.350 62.450 -23.150 ;
        RECT 54.850 -23.550 55.250 -23.350 ;
        RECT 62.050 -23.550 62.450 -23.350 ;
        RECT 39.650 -26.450 40.050 -23.900 ;
        RECT 42.550 -26.450 42.950 -23.800 ;
        RECT 45.450 -26.450 45.850 -23.800 ;
        RECT 49.750 -26.450 50.150 -23.900 ;
        RECT 54.050 -26.450 54.450 -23.900 ;
        RECT 56.950 -26.450 57.350 -23.800 ;
        RECT 59.850 -26.450 60.250 -23.800 ;
        RECT 64.150 -26.450 64.550 -23.900 ;
        RECT 68.200 -26.450 68.700 -3.850 ;
        RECT 80.970 -13.010 81.270 -12.160 ;
        RECT 96.150 -12.400 96.550 -12.250 ;
        RECT 97.800 -12.400 98.200 -12.350 ;
        RECT 84.310 -12.520 84.600 -12.475 ;
        RECT 86.410 -12.520 86.700 -12.475 ;
        RECT 87.980 -12.520 88.270 -12.475 ;
        RECT 84.310 -12.660 88.270 -12.520 ;
        RECT 84.310 -12.705 84.600 -12.660 ;
        RECT 86.410 -12.705 86.700 -12.660 ;
        RECT 87.980 -12.705 88.270 -12.660 ;
        RECT 96.150 -12.750 98.200 -12.400 ;
        RECT 80.000 -13.100 80.400 -13.050 ;
        RECT 77.400 -13.450 80.400 -13.100 ;
        RECT 80.980 -13.110 81.270 -13.010 ;
        RECT 84.705 -12.860 84.995 -12.815 ;
        RECT 85.895 -12.860 86.185 -12.815 ;
        RECT 88.415 -12.860 88.705 -12.815 ;
        RECT 84.705 -13.000 88.705 -12.860 ;
        RECT 84.705 -13.045 84.995 -13.000 ;
        RECT 85.895 -13.045 86.185 -13.000 ;
        RECT 88.415 -13.045 88.705 -13.000 ;
        RECT 80.980 -13.410 82.860 -13.110 ;
        RECT 77.400 -13.600 77.900 -13.450 ;
        RECT 80.000 -13.500 80.400 -13.450 ;
        RECT 82.630 -13.700 82.860 -13.410 ;
        RECT 85.090 -13.700 85.370 -13.410 ;
        RECT 95.350 -13.450 96.100 -13.100 ;
        RECT 95.350 -13.550 95.650 -13.450 ;
        RECT 82.630 -14.000 85.370 -13.700 ;
        RECT 93.600 -13.850 95.650 -13.550 ;
        RECT 39.650 -26.850 68.700 -26.450 ;
        RECT 34.200 -28.450 45.550 -28.050 ;
        RECT 45.150 -29.700 45.550 -28.450 ;
        RECT 45.150 -29.710 47.250 -29.700 ;
        RECT 45.150 -30.070 47.580 -29.710 ;
        RECT 48.200 -29.750 48.450 -28.750 ;
        RECT 49.850 -29.750 54.450 -29.600 ;
        RECT 48.200 -29.950 54.450 -29.750 ;
        RECT 48.285 -29.960 54.450 -29.950 ;
        RECT 45.150 -30.100 47.250 -30.070 ;
        RECT 49.850 -30.100 54.450 -29.960 ;
        RECT 53.950 -32.350 54.450 -30.100 ;
        RECT 60.060 -31.820 60.350 -31.775 ;
        RECT 62.160 -31.820 62.450 -31.775 ;
        RECT 63.730 -31.820 64.020 -31.775 ;
        RECT 60.060 -31.960 64.020 -31.820 ;
        RECT 60.060 -32.005 60.350 -31.960 ;
        RECT 62.160 -32.005 62.450 -31.960 ;
        RECT 63.730 -32.005 64.020 -31.960 ;
        RECT 60.455 -32.160 60.745 -32.115 ;
        RECT 61.645 -32.160 61.935 -32.115 ;
        RECT 64.165 -32.160 64.455 -32.115 ;
        RECT 60.455 -32.300 64.455 -32.160 ;
        RECT 60.455 -32.345 60.745 -32.300 ;
        RECT 61.645 -32.345 61.935 -32.300 ;
        RECT 64.165 -32.345 64.455 -32.300 ;
        RECT 52.200 -32.650 55.400 -32.350 ;
        RECT 33.950 -33.200 34.350 -32.700 ;
        RECT 34.650 -32.850 35.050 -32.750 ;
        RECT 36.450 -32.850 36.850 -32.750 ;
        RECT 34.650 -33.400 36.850 -32.850 ;
        RECT 34.650 -33.550 35.050 -33.400 ;
        RECT 36.450 -33.550 36.850 -33.400 ;
        RECT 26.300 -36.450 26.700 -33.550 ;
        RECT 30.050 -34.450 32.250 -33.950 ;
        RECT 30.050 -34.550 30.450 -34.450 ;
        RECT 31.850 -34.550 32.250 -34.450 ;
        RECT 35.550 -34.550 37.750 -33.950 ;
        RECT 39.450 -36.450 39.850 -32.750 ;
        RECT 40.150 -36.450 40.550 -33.600 ;
        RECT 52.200 -34.350 52.500 -32.650 ;
        RECT 55.000 -32.750 55.400 -32.650 ;
        RECT 60.750 -32.900 61.250 -32.550 ;
        RECT 58.100 -33.250 61.250 -32.900 ;
        RECT 58.100 -33.450 58.650 -33.250 ;
        RECT 66.400 -33.350 71.350 -32.850 ;
        RECT 52.200 -34.650 56.150 -34.350 ;
        RECT 26.300 -36.850 40.550 -36.450 ;
        RECT 55.850 -36.700 56.150 -34.650 ;
        RECT 68.500 -35.650 69.000 -34.500 ;
        RECT 64.950 -35.900 69.000 -35.650 ;
        RECT 58.660 -36.020 58.950 -35.975 ;
        RECT 60.760 -36.020 61.050 -35.975 ;
        RECT 62.330 -36.020 62.620 -35.975 ;
        RECT 58.660 -36.160 62.620 -36.020 ;
        RECT 58.660 -36.205 58.950 -36.160 ;
        RECT 60.760 -36.205 61.050 -36.160 ;
        RECT 62.330 -36.205 62.620 -36.160 ;
        RECT 58.150 -36.700 58.550 -36.350 ;
        RECT 59.055 -36.360 59.345 -36.315 ;
        RECT 60.245 -36.360 60.535 -36.315 ;
        RECT 62.765 -36.360 63.055 -36.315 ;
        RECT 59.055 -36.500 63.055 -36.360 ;
        RECT 59.055 -36.545 59.345 -36.500 ;
        RECT 60.245 -36.545 60.535 -36.500 ;
        RECT 62.765 -36.545 63.055 -36.500 ;
        RECT 55.850 -37.000 58.550 -36.700 ;
        RECT 59.450 -37.250 59.850 -36.650 ;
        RECT 57.100 -37.500 59.850 -37.250 ;
        RECT 64.950 -36.700 65.400 -35.900 ;
        RECT 64.950 -37.450 65.450 -36.700 ;
        RECT 28.550 -39.200 33.950 -38.700 ;
        RECT 25.050 -40.250 25.450 -39.750 ;
        RECT 25.750 -39.950 26.150 -39.800 ;
        RECT 27.550 -39.950 27.950 -39.800 ;
        RECT 25.750 -40.450 27.950 -39.950 ;
        RECT 25.750 -40.600 26.150 -40.450 ;
        RECT 27.550 -40.600 27.950 -40.450 ;
        RECT 19.300 -42.450 19.700 -40.950 ;
        RECT 25.750 -43.150 26.150 -43.000 ;
        RECT 27.550 -43.150 27.950 -43.000 ;
        RECT 25.750 -43.650 27.950 -43.150 ;
        RECT 25.750 -43.800 26.150 -43.650 ;
        RECT 27.550 -43.800 27.950 -43.650 ;
        RECT 28.550 -44.200 29.050 -39.200 ;
        RECT 30.550 -40.150 30.950 -39.950 ;
        RECT 32.350 -40.150 32.750 -39.950 ;
        RECT 30.550 -40.650 32.750 -40.150 ;
        RECT 30.550 -40.800 30.950 -40.650 ;
        RECT 32.350 -40.800 32.750 -40.650 ;
        RECT 33.450 -42.350 33.950 -39.200 ;
        RECT 57.100 -39.750 57.600 -37.500 ;
        RECT 68.000 -37.600 68.500 -37.200 ;
        RECT 70.850 -39.750 71.350 -33.350 ;
        RECT 34.400 -40.450 34.800 -39.950 ;
        RECT 36.200 -40.450 36.600 -39.950 ;
        RECT 38.900 -40.400 39.300 -39.900 ;
        RECT 39.600 -40.000 40.000 -39.850 ;
        RECT 41.400 -40.000 41.800 -39.850 ;
        RECT 34.400 -40.950 36.600 -40.450 ;
        RECT 39.600 -40.500 41.800 -40.000 ;
        RECT 57.100 -40.250 71.350 -39.750 ;
        RECT 39.600 -40.650 40.000 -40.500 ;
        RECT 41.400 -40.650 41.800 -40.500 ;
        RECT 34.400 -41.100 34.800 -40.950 ;
        RECT 36.200 -41.100 36.600 -40.950 ;
        RECT 72.300 -41.400 72.800 -34.500 ;
        RECT 82.130 -35.650 82.420 -35.605 ;
        RECT 83.990 -35.650 84.280 -35.605 ;
        RECT 86.770 -35.650 87.060 -35.605 ;
        RECT 82.130 -35.790 87.060 -35.650 ;
        RECT 82.130 -35.835 82.420 -35.790 ;
        RECT 83.990 -35.835 84.280 -35.790 ;
        RECT 86.770 -35.835 87.060 -35.790 ;
        RECT 94.100 -35.830 96.400 -35.480 ;
        RECT 74.200 -36.900 75.150 -36.000 ;
        RECT 80.600 -36.480 83.750 -36.080 ;
        RECT 86.770 -36.330 87.060 -36.285 ;
        RECT 84.525 -36.470 87.060 -36.330 ;
        RECT 53.800 -41.900 72.800 -41.400 ;
        RECT 79.300 -41.430 79.750 -41.380 ;
        RECT 78.900 -41.780 79.750 -41.430 ;
        RECT 79.300 -41.830 79.750 -41.780 ;
        RECT 30.950 -42.850 32.350 -42.350 ;
        RECT 33.450 -42.850 36.200 -42.350 ;
        RECT 39.600 -43.200 40.000 -43.050 ;
        RECT 41.400 -43.200 41.800 -43.050 ;
        RECT 39.600 -43.700 41.800 -43.200 ;
        RECT 39.600 -43.850 40.000 -43.700 ;
        RECT 41.400 -43.850 41.800 -43.700 ;
        RECT 53.800 -44.050 54.300 -41.900 ;
        RECT 80.600 -43.330 80.950 -36.480 ;
        RECT 84.525 -36.625 84.740 -36.470 ;
        RECT 86.770 -36.515 87.060 -36.470 ;
        RECT 82.590 -36.670 82.880 -36.625 ;
        RECT 84.450 -36.670 84.740 -36.625 ;
        RECT 85.370 -36.630 85.660 -36.625 ;
        RECT 82.590 -36.810 84.740 -36.670 ;
        RECT 82.590 -36.855 82.880 -36.810 ;
        RECT 84.450 -36.855 84.740 -36.810 ;
        RECT 85.300 -36.670 85.800 -36.630 ;
        RECT 88.630 -36.670 88.920 -36.625 ;
        RECT 85.300 -36.810 88.920 -36.670 ;
        RECT 85.300 -37.080 85.800 -36.810 ;
        RECT 88.630 -36.855 88.920 -36.810 ;
        RECT 92.050 -39.080 92.400 -36.230 ;
        RECT 84.700 -39.430 92.400 -39.080 ;
        RECT 84.700 -41.080 85.050 -39.430 ;
        RECT 84.700 -41.430 87.600 -41.080 ;
        RECT 86.650 -42.280 87.000 -41.930 ;
        RECT 87.250 -41.980 87.600 -41.430 ;
        RECT 91.900 -41.880 92.200 -41.180 ;
        RECT 93.500 -41.880 94.000 -41.800 ;
        RECT 87.150 -42.230 87.700 -41.980 ;
        RECT 91.900 -42.230 94.000 -41.880 ;
        RECT 91.900 -42.240 92.200 -42.230 ;
        RECT 60.060 -43.520 60.350 -43.475 ;
        RECT 62.160 -43.520 62.450 -43.475 ;
        RECT 63.730 -43.520 64.020 -43.475 ;
        RECT 60.060 -43.660 64.020 -43.520 ;
        RECT 60.060 -43.705 60.350 -43.660 ;
        RECT 62.160 -43.705 62.450 -43.660 ;
        RECT 63.730 -43.705 64.020 -43.660 ;
        RECT 77.950 -43.630 80.950 -43.330 ;
        RECT 84.700 -42.630 87.000 -42.280 ;
        RECT 93.500 -42.300 94.000 -42.230 ;
        RECT 60.455 -43.860 60.745 -43.815 ;
        RECT 61.645 -43.860 61.935 -43.815 ;
        RECT 64.165 -43.860 64.455 -43.815 ;
        RECT 60.455 -44.000 64.455 -43.860 ;
        RECT 60.455 -44.045 60.745 -44.000 ;
        RECT 61.645 -44.045 61.935 -44.000 ;
        RECT 64.165 -44.045 64.455 -44.000 ;
        RECT 26.150 -44.700 29.050 -44.200 ;
        RECT 40.000 -44.750 41.800 -44.250 ;
        RECT 19.700 -46.150 20.550 -45.800 ;
        RECT 26.450 -45.950 27.250 -45.250 ;
        RECT 19.700 -47.800 20.200 -46.150 ;
        RECT 26.650 -49.150 27.050 -45.950 ;
        RECT 41.400 -46.700 41.800 -44.750 ;
        RECT 52.200 -44.350 55.400 -44.050 ;
        RECT 52.200 -46.050 52.500 -44.350 ;
        RECT 55.000 -44.450 55.400 -44.350 ;
        RECT 60.750 -44.600 61.250 -44.250 ;
        RECT 58.100 -44.950 61.250 -44.600 ;
        RECT 58.100 -45.150 58.650 -44.950 ;
        RECT 66.400 -45.050 71.350 -44.550 ;
        RECT 52.200 -46.350 56.150 -46.050 ;
        RECT 55.850 -48.400 56.150 -46.350 ;
        RECT 68.500 -47.350 69.000 -46.200 ;
        RECT 64.950 -47.600 69.000 -47.350 ;
        RECT 58.660 -47.720 58.950 -47.675 ;
        RECT 60.760 -47.720 61.050 -47.675 ;
        RECT 62.330 -47.720 62.620 -47.675 ;
        RECT 58.660 -47.860 62.620 -47.720 ;
        RECT 58.660 -47.905 58.950 -47.860 ;
        RECT 60.760 -47.905 61.050 -47.860 ;
        RECT 62.330 -47.905 62.620 -47.860 ;
        RECT 58.150 -48.400 58.550 -48.050 ;
        RECT 59.055 -48.060 59.345 -48.015 ;
        RECT 60.245 -48.060 60.535 -48.015 ;
        RECT 62.765 -48.060 63.055 -48.015 ;
        RECT 59.055 -48.200 63.055 -48.060 ;
        RECT 59.055 -48.245 59.345 -48.200 ;
        RECT 60.245 -48.245 60.535 -48.200 ;
        RECT 62.765 -48.245 63.055 -48.200 ;
        RECT 55.850 -48.700 58.550 -48.400 ;
        RECT 59.450 -48.950 59.850 -48.350 ;
        RECT 26.650 -49.220 28.100 -49.150 ;
        RECT 57.100 -49.200 59.850 -48.950 ;
        RECT 64.950 -48.400 65.400 -47.600 ;
        RECT 64.950 -49.150 65.450 -48.400 ;
        RECT 26.650 -49.470 30.065 -49.220 ;
        RECT 26.650 -49.550 28.100 -49.470 ;
        RECT 57.100 -51.450 57.600 -49.200 ;
        RECT 68.000 -49.300 68.500 -48.900 ;
        RECT 70.850 -51.450 71.350 -45.050 ;
        RECT 77.950 -45.780 78.300 -43.630 ;
        RECT 84.700 -44.330 85.050 -42.630 ;
        RECT 96.050 -44.130 96.400 -35.830 ;
        RECT 80.950 -44.680 85.050 -44.330 ;
        RECT 91.700 -44.480 96.400 -44.130 ;
        RECT 80.950 -45.730 81.300 -44.680 ;
        RECT 77.950 -46.130 80.000 -45.780 ;
        RECT 80.950 -46.130 82.400 -45.730 ;
        RECT 83.940 -46.020 84.230 -45.975 ;
        RECT 87.200 -46.020 87.700 -45.680 ;
        RECT 83.940 -46.160 87.700 -46.020 ;
        RECT 83.940 -46.205 84.230 -46.160 ;
        RECT 87.200 -46.180 87.700 -46.160 ;
        RECT 88.120 -46.020 88.410 -45.975 ;
        RECT 89.980 -46.020 90.270 -45.975 ;
        RECT 88.120 -46.160 90.270 -46.020 ;
        RECT 87.200 -46.205 87.490 -46.180 ;
        RECT 88.120 -46.205 88.410 -46.160 ;
        RECT 89.980 -46.205 90.270 -46.160 ;
        RECT 85.800 -46.360 86.090 -46.315 ;
        RECT 88.120 -46.360 88.335 -46.205 ;
        RECT 85.800 -46.500 88.335 -46.360 ;
        RECT 85.800 -46.545 86.090 -46.500 ;
        RECT 89.100 -46.530 89.500 -46.330 ;
        RECT 91.700 -46.530 92.050 -44.480 ;
        RECT 108.050 -46.150 108.550 -12.400 ;
        RECT 89.100 -46.830 92.050 -46.530 ;
        RECT 92.400 -46.580 94.050 -46.230 ;
        RECT 89.100 -46.880 90.300 -46.830 ;
        RECT 90.900 -46.880 92.050 -46.830 ;
        RECT 85.800 -47.040 86.090 -46.995 ;
        RECT 88.580 -47.040 88.870 -46.995 ;
        RECT 90.440 -47.040 90.730 -46.995 ;
        RECT 85.800 -47.180 90.730 -47.040 ;
        RECT 85.800 -47.225 86.090 -47.180 ;
        RECT 88.580 -47.225 88.870 -47.180 ;
        RECT 90.440 -47.225 90.730 -47.180 ;
        RECT 93.700 -47.380 94.050 -46.580 ;
        RECT 95.400 -46.650 108.550 -46.150 ;
        RECT 57.100 -51.950 71.350 -51.450 ;
        RECT 108.050 -62.450 108.550 -46.650 ;
        RECT 2.350 -62.950 108.550 -62.450 ;
      LAYER met2 ;
        RECT -8.050 -15.130 -7.550 -14.580 ;
        RECT -8.050 -16.280 -7.700 -15.130 ;
        RECT -11.200 -16.630 -7.700 -16.280 ;
        RECT -14.050 -19.380 -13.600 -19.330 ;
        RECT -11.200 -19.380 -10.850 -16.630 ;
        RECT -14.050 -19.730 -10.850 -19.380 ;
        RECT -14.050 -19.780 -13.600 -19.730 ;
        RECT -11.200 -21.680 -10.850 -19.730 ;
        RECT -0.100 -20.200 5.000 -19.800 ;
        RECT -11.200 -22.030 -5.800 -21.680 ;
        RECT -6.150 -23.630 -5.800 -22.030 ;
        RECT -6.150 -24.130 -5.650 -23.630 ;
        RECT 4.600 -38.350 5.000 -20.200 ;
        RECT 77.400 -31.500 77.900 -13.100 ;
        RECT 77.400 -32.000 98.500 -31.500 ;
        RECT 68.500 -35.000 72.800 -34.500 ;
        RECT 74.200 -36.900 75.150 -36.000 ;
        RECT 4.600 -38.750 19.700 -38.350 ;
        RECT 19.300 -40.900 19.700 -38.750 ;
        RECT 19.250 -41.350 19.750 -40.900 ;
        RECT 74.345 -46.200 74.860 -36.900 ;
        RECT 85.300 -37.180 85.800 -36.630 ;
        RECT 85.300 -38.330 85.650 -37.180 ;
        RECT 82.150 -38.680 85.650 -38.330 ;
        RECT 79.300 -41.430 79.750 -41.380 ;
        RECT 82.150 -41.430 82.500 -38.680 ;
        RECT 79.300 -41.780 82.500 -41.430 ;
        RECT 79.300 -41.830 79.750 -41.780 ;
        RECT 82.150 -43.730 82.500 -41.780 ;
        RECT 98.000 -41.800 98.500 -32.000 ;
        RECT 93.500 -42.300 98.500 -41.800 ;
        RECT 82.150 -44.080 87.550 -43.730 ;
        RECT 87.200 -45.680 87.550 -44.080 ;
        RECT 87.200 -46.180 87.700 -45.680 ;
        RECT 68.500 -46.700 74.860 -46.200 ;
        RECT 74.345 -46.705 74.860 -46.700 ;
  END
END system
END LIBRARY

