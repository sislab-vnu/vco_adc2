magic
tech sky130A
magscale 1 2
timestamp 1730705417
<< locali >>
rect -2830 4030 3060 4050
rect -2830 3970 -2810 4030
rect -2750 3970 -2710 4030
rect -2650 3970 2740 4030
rect 2800 3970 2860 4030
rect 2920 3970 2980 4030
rect 3040 3970 3060 4030
rect -2830 3950 3060 3970
rect -2830 3930 -2730 3950
rect -2830 3870 -2810 3930
rect -2750 3870 -2730 3930
rect -2830 3850 -2730 3870
rect 2320 930 2420 3950
rect 2320 830 6030 930
rect 5930 -1180 6030 830
rect 5930 -1280 7040 -1180
rect 1130 -1560 6110 -1540
rect 1130 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 1130 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 6030 -1700 6110 -1680
rect 6940 -1690 7040 -1280
rect 6940 -1710 8290 -1690
rect 6940 -1770 8010 -1710
rect 8070 -1770 8110 -1710
rect 8170 -1770 8210 -1710
rect 8270 -1770 8290 -1710
rect 6940 -1790 8290 -1770
rect 1470 -2150 2740 -2130
rect 1470 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 1470 -2220 2740 -2210
rect 1530 -2230 2740 -2220
rect 1580 -2420 3950 -2400
rect 1580 -2480 3770 -2420
rect 3830 -2480 3870 -2420
rect 3930 -2480 3950 -2420
rect 1580 -2500 3950 -2480
rect 3850 -2520 3950 -2500
rect 3850 -2580 3870 -2520
rect 3930 -2580 3950 -2520
rect 3850 -2600 3950 -2580
rect 3850 -4790 3950 -4770
rect 3850 -4850 3870 -4790
rect 3930 -4850 3950 -4790
rect 3850 -4870 3950 -4850
rect 2080 -4890 3950 -4870
rect 2080 -4950 2100 -4890
rect 2160 -4950 2220 -4890
rect 2280 -4950 2340 -4890
rect 2400 -4950 3870 -4890
rect 3930 -4950 3950 -4890
rect 2080 -4970 3950 -4950
rect 3850 -4990 3950 -4970
rect 3850 -5050 3870 -4990
rect 3930 -5050 3950 -4990
rect 860 -5680 1060 -5050
rect 3850 -5070 3950 -5050
rect 860 -5720 880 -5680
rect 920 -5720 1000 -5680
rect 1040 -5720 1060 -5680
rect 860 -5810 1060 -5720
rect 860 -5850 880 -5810
rect 920 -5850 1000 -5810
rect 1040 -5850 1060 -5810
rect 860 -5870 1060 -5850
rect -2240 -6750 -1830 -6740
rect -2240 -6760 -1820 -6750
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -1820 -6760
rect -2240 -6820 -1820 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -2240 -6900 -2160 -6880
rect -2830 -7690 -2730 -7670
rect -2830 -7750 -2810 -7690
rect -2750 -7750 -2730 -7690
rect -2830 -7770 -2730 -7750
rect -2830 -7790 -1890 -7770
rect -2830 -7850 -2810 -7790
rect -2750 -7850 -2710 -7790
rect -2650 -7850 -2070 -7790
rect -2010 -7850 -1970 -7790
rect -1910 -7850 -1890 -7790
rect -2830 -7870 -1890 -7850
rect 1260 -7890 2370 -7870
rect 1260 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 1260 -7950 2370 -7930
rect 16280 -7900 17170 -7870
rect 16280 -7940 16310 -7900
rect 16350 -7940 16390 -7900
rect 16430 -7940 17170 -7900
rect 16280 -7970 17170 -7940
rect 16280 -7980 16380 -7970
rect 16280 -8020 16310 -7980
rect 16350 -8020 16380 -7980
rect 16280 -8050 16380 -8020
rect 3850 -8650 3950 -8630
rect 3850 -8710 3870 -8650
rect 3930 -8710 3950 -8650
rect 3850 -8730 3950 -8710
rect 1580 -8750 3950 -8730
rect 1580 -8810 3770 -8750
rect 3830 -8810 3870 -8750
rect 3930 -8810 3950 -8750
rect 1580 -8830 3950 -8810
rect 17070 -9960 17170 -7970
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect 17000 -10040 17170 -10020
rect 17000 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect 17000 -10100 17170 -10080
<< viali >>
rect -1090 8010 -1050 8050
rect -1010 8010 -970 8050
rect -930 8010 -890 8050
rect -850 8010 -810 8050
rect -770 8010 -730 8050
rect 3040 8010 3080 8050
rect 3120 8010 3160 8050
rect 3200 8010 3240 8050
rect 3280 8010 3320 8050
rect 3360 8010 3400 8050
rect 11060 8010 11100 8050
rect 11140 8010 11180 8050
rect 11220 8010 11260 8050
rect 11300 8010 11340 8050
rect 11380 8010 11420 8050
rect 15890 8010 15930 8050
rect 15970 8010 16010 8050
rect 16050 8010 16090 8050
rect 16130 8010 16170 8050
rect 16210 8010 16250 8050
rect -2810 3970 -2750 4030
rect -2710 3970 -2650 4030
rect 2740 3970 2800 4030
rect 2860 3970 2920 4030
rect 2980 3970 3040 4030
rect -2810 3870 -2750 3930
rect -2000 -470 -1960 -430
rect -1920 -470 -1880 -430
rect 1150 -1600 1190 -1560
rect 1230 -1600 1270 -1560
rect 5970 -1600 6010 -1560
rect 6050 -1600 6090 -1560
rect 6050 -1680 6090 -1640
rect 8010 -1770 8070 -1710
rect 8110 -1770 8170 -1710
rect 8210 -1770 8270 -1710
rect 2420 -2210 2480 -2150
rect 2540 -2210 2600 -2150
rect 2660 -2210 2720 -2150
rect 3770 -2480 3830 -2420
rect 3870 -2480 3930 -2420
rect 3870 -2580 3930 -2520
rect 3870 -4850 3930 -4790
rect 2100 -4950 2160 -4890
rect 2220 -4950 2280 -4890
rect 2340 -4950 2400 -4890
rect 3870 -4950 3930 -4890
rect 3870 -5050 3930 -4990
rect 880 -5720 920 -5680
rect 1000 -5720 1040 -5680
rect 880 -5850 920 -5810
rect 1000 -5850 1040 -5810
rect -2220 -6800 -2180 -6760
rect -2140 -6800 -2100 -6760
rect -2220 -6880 -2180 -6840
rect -2810 -7750 -2750 -7690
rect -2810 -7850 -2750 -7790
rect -2710 -7850 -2650 -7790
rect -2070 -7850 -2010 -7790
rect -1970 -7850 -1910 -7790
rect 1280 -7930 1320 -7890
rect 1360 -7930 1400 -7890
rect 1440 -7930 1480 -7890
rect 2150 -7930 2190 -7890
rect 2230 -7930 2270 -7890
rect 2310 -7930 2350 -7890
rect 16310 -7940 16350 -7900
rect 16390 -7940 16430 -7900
rect 16310 -8020 16350 -7980
rect 3870 -8710 3930 -8650
rect 3770 -8810 3830 -8750
rect 3870 -8810 3930 -8750
rect 17100 -10000 17140 -9960
rect 17020 -10080 17060 -10040
rect 17100 -10080 17140 -10040
<< metal1 >>
rect -1110 8060 -710 8070
rect -1110 8000 -1100 8060
rect -1040 8050 -980 8060
rect -920 8050 -860 8060
rect -800 8050 -710 8060
rect -1040 8010 -1010 8050
rect -890 8010 -860 8050
rect -800 8010 -770 8050
rect -730 8010 -710 8050
rect -1040 8000 -980 8010
rect -920 8000 -860 8010
rect -800 8000 -710 8010
rect -1110 7990 -710 8000
rect 3020 8060 3420 8070
rect 3020 8000 3030 8060
rect 3090 8050 3190 8060
rect 3250 8050 3350 8060
rect 3090 8010 3120 8050
rect 3160 8010 3190 8050
rect 3250 8010 3280 8050
rect 3320 8010 3350 8050
rect 3090 8000 3190 8010
rect 3250 8000 3350 8010
rect 3410 8000 3420 8060
rect 3020 7990 3420 8000
rect 11040 8060 11440 8070
rect 11040 8000 11050 8060
rect 11110 8050 11210 8060
rect 11270 8050 11370 8060
rect 11110 8010 11140 8050
rect 11180 8010 11210 8050
rect 11270 8010 11300 8050
rect 11340 8010 11370 8050
rect 11110 8000 11210 8010
rect 11270 8000 11370 8010
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8060 16270 8070
rect 15870 8000 15880 8060
rect 15940 8050 16040 8060
rect 16100 8050 16200 8060
rect 15940 8010 15970 8050
rect 16010 8010 16040 8050
rect 16100 8010 16130 8050
rect 16170 8010 16200 8050
rect 15940 8000 16040 8010
rect 16100 8000 16200 8010
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 6900 4980 7140 5000
rect 6900 4920 6920 4980
rect 6980 4920 7040 4980
rect 7100 4920 7140 4980
rect 6900 4880 7140 4920
rect 6900 4820 6920 4880
rect 6980 4820 7040 4880
rect 7100 4820 7140 4880
rect 6900 4800 7140 4820
rect -2830 4030 -2630 4050
rect -2830 3970 -2810 4030
rect -2750 3970 -2710 4030
rect -2650 3970 -2630 4030
rect -2830 3930 -2630 3970
rect 2710 4030 3060 4050
rect 2710 3970 2740 4030
rect 2800 3970 2860 4030
rect 2920 3970 2980 4030
rect 3040 3970 3060 4030
rect 2710 3950 3060 3970
rect -2830 3870 -2810 3930
rect -2750 3870 -2630 3930
rect -2830 3770 -2630 3870
rect -2830 3670 -2790 3770
rect -2690 3670 -2630 3770
rect -2830 3570 -2630 3670
rect -2830 3470 -2790 3570
rect -2690 3470 -2630 3570
rect -2830 3370 -2630 3470
rect -2830 3270 -2790 3370
rect -2690 3270 -2630 3370
rect -2830 -1430 -2630 3270
rect -2020 -410 -1920 2100
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 -130 -1080 1010
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 -120 80 1000
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 -130 1290 1020
rect -2020 -430 -1860 -410
rect -2020 -470 -2000 -430
rect -1960 -470 -1920 -430
rect -1880 -470 -1860 -430
rect -2020 -490 -1860 -470
rect -2830 -1456 -2000 -1430
rect -2830 -1526 -1875 -1456
rect -2830 -1530 -2000 -1526
rect -2830 -7690 -2630 -1530
rect 970 -1560 1290 -1540
rect 970 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 1290 -1560
rect 970 -1620 1290 -1600
rect 5950 -1560 6110 -1540
rect 5950 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 5950 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 2400 -2150 2740 -2130
rect 2400 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 2400 -2230 2740 -2210
rect 2360 -3100 2760 -2230
rect 3750 -2420 3950 -2400
rect 3750 -2480 3770 -2420
rect 3830 -2480 3870 -2420
rect 3930 -2480 3950 -2420
rect 3750 -2500 3950 -2480
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3480 2760 -3280
rect 3850 -2520 3950 -2500
rect 3850 -2580 3870 -2520
rect 3930 -2580 3950 -2520
rect -2320 -4490 -1920 -3900
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4800 -1920 -4550
rect -1770 -4210 -1570 -4190
rect -1770 -4310 -1730 -4210
rect -1630 -4310 -1570 -4210
rect -1770 -4380 -1570 -4310
rect -1770 -4480 -1730 -4380
rect -1630 -4480 -1570 -4380
rect -1770 -4540 -1570 -4480
rect -1770 -4640 -1730 -4540
rect -1630 -4640 -1570 -4540
rect -1770 -4660 -1570 -4640
rect 3850 -4790 3950 -2580
rect 3850 -4850 3870 -4790
rect 3930 -4850 3950 -4790
rect 2080 -4890 2420 -4870
rect 2080 -4950 2100 -4890
rect 2160 -4950 2220 -4890
rect 2280 -4950 2340 -4890
rect 2400 -4950 2420 -4890
rect 2080 -4970 2420 -4950
rect 3850 -4890 3950 -4850
rect 3850 -4950 3870 -4890
rect 3930 -4950 3950 -4890
rect 6030 -4830 6110 -1680
rect 7990 -1710 8290 -1690
rect 7990 -1770 8010 -1710
rect 8070 -1770 8110 -1710
rect 8170 -1770 8210 -1710
rect 8270 -1770 8290 -1710
rect 7990 -1790 8290 -1770
rect 13160 -3580 13250 -3540
rect 13160 -3640 13170 -3580
rect 13230 -3640 13250 -3580
rect 13160 -3700 13250 -3640
rect 13160 -3760 13170 -3700
rect 13230 -3760 13250 -3700
rect 13160 -3890 13250 -3760
rect 6540 -4480 6740 -4460
rect 6540 -4540 6560 -4480
rect 6620 -4540 6660 -4480
rect 6720 -4500 6740 -4480
rect 6720 -4540 8190 -4500
rect 6540 -4580 8190 -4540
rect 6540 -4640 6560 -4580
rect 6620 -4640 6660 -4580
rect 6720 -4600 8190 -4580
rect 6720 -4640 6740 -4600
rect 6540 -4660 6740 -4640
rect 6030 -4910 6520 -4830
rect 3850 -4990 3950 -4950
rect -1790 -6070 -1710 -5020
rect 3850 -5050 3870 -4990
rect 3930 -5050 3950 -4990
rect -1480 -5500 -1080 -5340
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5580 -1080 -5560
rect -90 -5500 310 -5340
rect -90 -5560 -60 -5500
rect 0 -5560 60 -5500
rect 120 -5560 180 -5500
rect 240 -5560 310 -5500
rect -90 -5580 310 -5560
rect 860 -5680 1280 -5670
rect 860 -5720 880 -5680
rect 920 -5720 1000 -5680
rect 1040 -5690 1280 -5680
rect 1040 -5720 1080 -5690
rect 860 -5750 1080 -5720
rect 1140 -5750 1200 -5690
rect 1260 -5750 1280 -5690
rect 860 -5790 1280 -5750
rect 860 -5810 1080 -5790
rect 860 -5850 880 -5810
rect 920 -5850 1000 -5810
rect 1040 -5850 1080 -5810
rect 1140 -5850 1200 -5790
rect 1260 -5850 1280 -5790
rect 860 -5870 1280 -5850
rect -1790 -6150 2370 -6070
rect -2830 -7750 -2810 -7690
rect -2750 -7750 -2630 -7690
rect -2830 -7790 -2630 -7750
rect -2830 -7850 -2810 -7790
rect -2750 -7850 -2710 -7790
rect -2650 -7850 -2630 -7790
rect -2830 -7870 -2630 -7850
rect -2240 -6760 -2080 -6740
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -2080 -6760
rect -2240 -6820 -2080 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -2240 -10020 -2160 -6880
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7170 -1480 -7150
rect -2100 -7790 -1890 -7770
rect -2100 -7850 -2070 -7790
rect -2010 -7850 -1970 -7790
rect -1910 -7850 -1890 -7790
rect -2100 -7870 -1890 -7850
rect 2290 -7870 2370 -6150
rect 970 -7890 1500 -7870
rect 970 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 1500 -7890
rect 970 -7950 1500 -7930
rect 2130 -7890 2370 -7870
rect 2130 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 2130 -7950 2370 -7930
rect 3850 -8650 3950 -5050
rect 6440 -7010 6520 -4910
rect 9100 -4950 9300 -4930
rect 9100 -5010 9120 -4950
rect 9180 -5010 9220 -4950
rect 9280 -5010 9300 -4950
rect 9100 -5050 9300 -5010
rect 9100 -5110 9120 -5050
rect 9180 -5110 9220 -5050
rect 9280 -5110 9300 -5050
rect 9100 -5130 9300 -5110
rect 16280 -7900 16490 -7870
rect 16280 -7940 16310 -7900
rect 16350 -7940 16390 -7900
rect 16430 -7940 16490 -7900
rect 16280 -7970 16490 -7940
rect 16280 -7980 16380 -7970
rect 16280 -8020 16310 -7980
rect 16350 -8020 16380 -7980
rect 16280 -8050 16380 -8020
rect 12250 -8140 12650 -8120
rect 12250 -8200 12280 -8140
rect 12340 -8200 12400 -8140
rect 12460 -8200 12520 -8140
rect 12580 -8200 12650 -8140
rect 12250 -8220 12650 -8200
rect 3850 -8710 3870 -8650
rect 3930 -8710 3950 -8650
rect 3850 -8730 3950 -8710
rect 3750 -8750 3950 -8730
rect 3750 -8810 3770 -8750
rect 3830 -8810 3870 -8750
rect 3930 -8810 3950 -8750
rect 3750 -8830 3950 -8810
rect -1640 -9170 -1240 -9050
rect -1640 -9230 -1610 -9170
rect -1550 -9230 -1490 -9170
rect -1430 -9230 -1370 -9170
rect -1310 -9230 -1240 -9170
rect -1640 -9370 -1240 -9230
rect 580 -9160 980 -9060
rect 580 -9220 610 -9160
rect 670 -9220 730 -9160
rect 790 -9220 850 -9160
rect 910 -9220 980 -9160
rect 580 -9250 980 -9220
rect 17070 -9960 17170 -9940
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect -2240 -10040 17170 -10020
rect -2240 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect -2240 -10100 17170 -10080
<< via1 >>
rect -1100 8050 -1040 8060
rect -980 8050 -920 8060
rect -860 8050 -800 8060
rect -1100 8010 -1090 8050
rect -1090 8010 -1050 8050
rect -1050 8010 -1040 8050
rect -980 8010 -970 8050
rect -970 8010 -930 8050
rect -930 8010 -920 8050
rect -860 8010 -850 8050
rect -850 8010 -810 8050
rect -810 8010 -800 8050
rect -1100 8000 -1040 8010
rect -980 8000 -920 8010
rect -860 8000 -800 8010
rect 3030 8050 3090 8060
rect 3190 8050 3250 8060
rect 3350 8050 3410 8060
rect 3030 8010 3040 8050
rect 3040 8010 3080 8050
rect 3080 8010 3090 8050
rect 3190 8010 3200 8050
rect 3200 8010 3240 8050
rect 3240 8010 3250 8050
rect 3350 8010 3360 8050
rect 3360 8010 3400 8050
rect 3400 8010 3410 8050
rect 3030 8000 3090 8010
rect 3190 8000 3250 8010
rect 3350 8000 3410 8010
rect 11050 8050 11110 8060
rect 11210 8050 11270 8060
rect 11370 8050 11430 8060
rect 11050 8010 11060 8050
rect 11060 8010 11100 8050
rect 11100 8010 11110 8050
rect 11210 8010 11220 8050
rect 11220 8010 11260 8050
rect 11260 8010 11270 8050
rect 11370 8010 11380 8050
rect 11380 8010 11420 8050
rect 11420 8010 11430 8050
rect 11050 8000 11110 8010
rect 11210 8000 11270 8010
rect 11370 8000 11430 8010
rect 15880 8050 15940 8060
rect 16040 8050 16100 8060
rect 16200 8050 16260 8060
rect 15880 8010 15890 8050
rect 15890 8010 15930 8050
rect 15930 8010 15940 8050
rect 16040 8010 16050 8050
rect 16050 8010 16090 8050
rect 16090 8010 16100 8050
rect 16200 8010 16210 8050
rect 16210 8010 16250 8050
rect 16250 8010 16260 8050
rect 15880 8000 15940 8010
rect 16040 8000 16100 8010
rect 16200 8000 16260 8010
rect 6920 4920 6980 4980
rect 7040 4920 7100 4980
rect 6920 4820 6980 4880
rect 7040 4820 7100 4880
rect 14700 4500 14760 4560
rect 14700 4380 14760 4440
rect 14700 4260 14760 4320
rect -2790 3670 -2690 3770
rect -2790 3470 -2690 3570
rect -2790 3270 -2690 3370
rect -1430 1010 -1360 1080
rect -1200 1010 -1130 1080
rect -270 1000 -200 1070
rect -50 1000 20 1070
rect 930 1020 990 1080
rect 1180 1020 1240 1080
rect 2390 -3160 2450 -3100
rect 2510 -3160 2570 -3100
rect 2630 -3160 2690 -3100
rect 2390 -3280 2450 -3220
rect 2510 -3280 2570 -3220
rect 2630 -3280 2690 -3220
rect -2280 -4550 -2220 -4490
rect -2030 -4550 -1970 -4490
rect -1730 -4310 -1630 -4210
rect -1730 -4480 -1630 -4380
rect -1730 -4640 -1630 -4540
rect 18530 -2080 18590 -2020
rect 18530 -2200 18590 -2140
rect 18530 -2320 18590 -2260
rect 13170 -3640 13230 -3580
rect 13170 -3760 13230 -3700
rect 6560 -4540 6620 -4480
rect 6660 -4540 6720 -4480
rect 6560 -4640 6620 -4580
rect 6660 -4640 6720 -4580
rect -1450 -5560 -1390 -5500
rect -1330 -5560 -1270 -5500
rect -1210 -5560 -1150 -5500
rect -60 -5560 0 -5500
rect 60 -5560 120 -5500
rect 180 -5560 240 -5500
rect 1080 -5750 1140 -5690
rect 1200 -5750 1260 -5690
rect 1080 -5850 1140 -5790
rect 1200 -5850 1260 -5790
rect -1930 -7150 -1870 -7090
rect -1810 -7150 -1750 -7090
rect -1690 -7150 -1630 -7090
rect -1570 -7150 -1510 -7090
rect 9120 -5010 9180 -4950
rect 9220 -5010 9280 -4950
rect 9120 -5110 9180 -5050
rect 9220 -5110 9280 -5050
rect 18530 -7070 18590 -7010
rect 18530 -7190 18590 -7130
rect 18530 -7310 18590 -7250
rect 12280 -8200 12340 -8140
rect 12400 -8200 12460 -8140
rect 12520 -8200 12580 -8140
rect -1610 -9230 -1550 -9170
rect -1490 -9230 -1430 -9170
rect -1370 -9230 -1310 -9170
rect 610 -9220 670 -9160
rect 730 -9220 790 -9160
rect 850 -9220 910 -9160
rect 8030 -9640 8090 -9580
rect 8150 -9640 8210 -9580
rect 8270 -9640 8330 -9580
rect 16090 -9640 16150 -9580
rect 16210 -9640 16270 -9580
rect 16330 -9640 16390 -9580
<< metal2 >>
rect 17342 35320 17710 36938
rect 17342 34920 22770 35320
rect 17342 34914 17710 34920
rect -1110 8180 -710 8210
rect -1110 8100 -1070 8180
rect -990 8100 -830 8180
rect -750 8100 -710 8180
rect -1110 8060 -710 8100
rect -1110 8000 -1100 8060
rect -1040 8000 -980 8060
rect -920 8000 -860 8060
rect -800 8000 -710 8060
rect -1110 7990 -710 8000
rect 3020 8190 3420 8210
rect 3020 8110 3060 8190
rect 3140 8110 3280 8190
rect 3360 8110 3420 8190
rect 3020 8060 3420 8110
rect 3020 8000 3030 8060
rect 3090 8000 3190 8060
rect 3250 8000 3350 8060
rect 3410 8000 3420 8060
rect 3020 7990 3420 8000
rect 11040 8190 11440 8220
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8060 11440 8110
rect 11040 8000 11050 8060
rect 11110 8000 11210 8060
rect 11270 8000 11370 8060
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8180 16270 8210
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8060 16270 8100
rect 15870 8000 15880 8060
rect 15940 8000 16040 8060
rect 16100 8000 16200 8060
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 22370 5000 22770 34920
rect 6900 4980 22770 5000
rect 6900 4920 6920 4980
rect 6980 4920 7040 4980
rect 7100 4920 22770 4980
rect 6900 4880 22770 4920
rect 6900 4820 6920 4880
rect 6980 4820 7040 4880
rect 7100 4820 22770 4880
rect 6900 4800 22770 4820
rect 14680 4570 14990 4630
rect 14680 4560 14830 4570
rect 14680 4500 14700 4560
rect 14760 4500 14830 4560
rect 14680 4470 14830 4500
rect 14930 4470 14990 4570
rect 14680 4440 14990 4470
rect 14680 4380 14700 4440
rect 14760 4380 14990 4440
rect 14680 4370 14990 4380
rect 14680 4320 14830 4370
rect 14680 4260 14700 4320
rect 14760 4270 14830 4320
rect 14930 4270 14990 4370
rect 14760 4260 14990 4270
rect 14680 4230 14990 4260
rect -7520 3770 -2630 3850
rect -7520 3670 -2790 3770
rect -2690 3670 -2630 3770
rect -7520 3570 -2630 3670
rect -7520 3470 -2790 3570
rect -2690 3470 -2630 3570
rect -7520 3450 -2630 3470
rect -7520 -16330 -7120 3450
rect -2830 3370 -2630 3450
rect -2830 3270 -2790 3370
rect -2690 3270 -2630 3370
rect -2830 3250 -2630 3270
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 960 -1080 1010
rect -1480 880 -1430 960
rect -1350 880 -1220 960
rect -1140 880 -1080 960
rect -1480 820 -1080 880
rect -1480 740 -1430 820
rect -1350 740 -1220 820
rect -1140 740 -1080 820
rect -1480 710 -1080 740
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 950 80 1000
rect -320 870 -270 950
rect -190 870 -50 950
rect 30 870 80 950
rect -320 810 80 870
rect -320 730 -270 810
rect -190 730 -50 810
rect 30 730 80 810
rect -320 710 80 730
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 980 1290 1020
rect 890 900 930 980
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 890 820 1290 900
rect 890 740 930 820
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 890 710 1290 740
rect 18510 -2000 18790 -1950
rect 18510 -2020 18650 -2000
rect 18510 -2080 18530 -2020
rect 18590 -2080 18650 -2020
rect 18730 -2080 18790 -2000
rect 18510 -2140 18790 -2080
rect 18510 -2200 18530 -2140
rect 18590 -2160 18790 -2140
rect 18590 -2200 18650 -2160
rect 18510 -2240 18650 -2200
rect 18730 -2240 18790 -2160
rect 18510 -2260 18790 -2240
rect 18510 -2320 18530 -2260
rect 18590 -2320 18790 -2260
rect 18510 -2350 18790 -2320
rect 2360 -3100 2760 -3080
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3340 2760 -3280
rect 2360 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect 2360 -3480 2760 -3420
rect -5170 -3760 -1570 -3560
rect -5170 -16330 -4770 -3760
rect -2320 -4220 -1920 -4190
rect -2320 -4300 -2290 -4220
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -2320 -4370 -1920 -4300
rect -2320 -4450 -2290 -4370
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -2320 -4490 -1920 -4450
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4590 -1920 -4550
rect -1770 -4210 -1570 -3760
rect 13160 -3570 13420 -3540
rect 13160 -3580 13300 -3570
rect 13160 -3640 13170 -3580
rect 13230 -3640 13300 -3580
rect 13160 -3650 13300 -3640
rect 13380 -3650 13420 -3570
rect 13160 -3700 13420 -3650
rect 13160 -3760 13170 -3700
rect 13230 -3760 13420 -3700
rect 13160 -3810 13420 -3760
rect 13160 -3890 13300 -3810
rect 13380 -3890 13420 -3810
rect 13160 -3940 13420 -3890
rect -1770 -4310 -1730 -4210
rect -1630 -4310 -1570 -4210
rect -1770 -4380 -1570 -4310
rect -1770 -4480 -1730 -4380
rect -1630 -4480 -1570 -4380
rect -1770 -4540 -1570 -4480
rect -1770 -4640 -1730 -4540
rect -1630 -4640 -1570 -4540
rect -1770 -4660 -1570 -4640
rect 4530 -4480 6740 -4460
rect 4530 -4540 6560 -4480
rect 6620 -4540 6660 -4480
rect 6720 -4540 6740 -4480
rect 4530 -4580 6740 -4540
rect 4530 -4640 6560 -4580
rect 6620 -4640 6660 -4580
rect 6720 -4640 6740 -4580
rect 4530 -4660 6740 -4640
rect -1480 -5500 -1080 -5470
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5630 -1080 -5560
rect -1480 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 -1080 -5630
rect -1480 -5770 -1080 -5710
rect -1480 -5850 -1430 -5770
rect -1350 -5850 -1230 -5770
rect -1150 -5850 -1080 -5770
rect -1480 -5870 -1080 -5850
rect -90 -5500 310 -5470
rect -90 -5560 -60 -5500
rect 0 -5560 60 -5500
rect 120 -5560 180 -5500
rect 240 -5560 310 -5500
rect -90 -5630 310 -5560
rect -90 -5710 -40 -5630
rect 40 -5710 160 -5630
rect 240 -5710 310 -5630
rect -90 -5770 310 -5710
rect -90 -5850 -40 -5770
rect 40 -5850 160 -5770
rect 240 -5850 310 -5770
rect -90 -5870 310 -5850
rect 1060 -5690 3230 -5670
rect 1060 -5750 1080 -5690
rect 1140 -5750 1200 -5690
rect 1260 -5750 3230 -5690
rect 1060 -5790 3230 -5750
rect 1060 -5850 1080 -5790
rect 1140 -5850 1200 -5790
rect 1260 -5850 3230 -5790
rect 1060 -5870 3230 -5850
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7210 -1480 -7150
rect -1960 -7290 -1930 -7210
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -1960 -7320 -1480 -7290
rect -1640 -9170 -1240 -9150
rect -1640 -9230 -1610 -9170
rect -1550 -9230 -1490 -9170
rect -1430 -9230 -1370 -9170
rect -1310 -9230 -1240 -9170
rect -1640 -9260 -1240 -9230
rect -1640 -9340 -1610 -9260
rect -1530 -9340 -1380 -9260
rect -1300 -9340 -1240 -9260
rect -1640 -9370 -1240 -9340
rect 580 -9160 980 -9140
rect 580 -9220 610 -9160
rect 670 -9220 730 -9160
rect 790 -9220 850 -9160
rect 910 -9220 980 -9160
rect 580 -9260 980 -9220
rect 580 -9340 610 -9260
rect 690 -9340 840 -9260
rect 920 -9340 980 -9260
rect 580 -9360 980 -9340
rect 2830 -16330 3230 -5870
rect -7590 -17526 -7038 -16330
rect -5198 -17526 -4646 -16330
rect 2806 -17526 3358 -16330
rect 4530 -63620 4930 -4660
rect 9100 -4890 11680 -4690
rect 9100 -4950 9300 -4890
rect 9100 -5010 9120 -4950
rect 9180 -5010 9220 -4950
rect 9280 -5010 9300 -4950
rect 9100 -5050 9300 -5010
rect 9100 -5110 9120 -5050
rect 9180 -5110 9220 -5050
rect 9280 -5110 9300 -5050
rect 9100 -5130 9300 -5110
rect 8000 -9580 8390 -9560
rect 8000 -9640 8030 -9580
rect 8090 -9640 8150 -9580
rect 8210 -9640 8270 -9580
rect 8330 -9640 8390 -9580
rect 8000 -9690 8390 -9640
rect 8000 -9770 8040 -9690
rect 8120 -9770 8260 -9690
rect 8340 -9770 8390 -9690
rect 8000 -9800 8390 -9770
rect 11480 -10560 11680 -4890
rect 18510 -7010 18760 -6940
rect 18510 -7070 18530 -7010
rect 18590 -7070 18760 -7010
rect 18510 -7130 18650 -7070
rect 18510 -7190 18530 -7130
rect 18590 -7150 18650 -7130
rect 18730 -7150 18760 -7070
rect 18590 -7190 18760 -7150
rect 18510 -7230 18760 -7190
rect 18510 -7250 18650 -7230
rect 18510 -7310 18530 -7250
rect 18590 -7310 18650 -7250
rect 18730 -7310 18760 -7230
rect 18510 -7340 18760 -7310
rect 12250 -8140 12650 -8120
rect 12250 -8200 12280 -8140
rect 12340 -8200 12400 -8140
rect 12460 -8200 12520 -8140
rect 12580 -8200 12650 -8140
rect 12250 -8230 12650 -8200
rect 12250 -8310 12270 -8230
rect 12350 -8310 12510 -8230
rect 12590 -8310 12650 -8230
rect 12250 -8320 12650 -8310
rect 16070 -9580 16460 -9560
rect 16070 -9640 16090 -9580
rect 16150 -9640 16210 -9580
rect 16270 -9640 16330 -9580
rect 16390 -9640 16460 -9580
rect 16070 -9690 16460 -9640
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9800 16460 -9770
rect 11480 -10650 26770 -10560
rect 11480 -10850 25420 -10650
rect 25620 -10850 25820 -10650
rect 26020 -10850 26220 -10650
rect 26420 -10850 26770 -10650
rect 11480 -10970 26770 -10850
rect 4530 -63720 26670 -63620
rect 4530 -63920 25350 -63720
rect 25550 -63920 25750 -63720
rect 25950 -63920 26150 -63720
rect 26350 -63920 26670 -63720
rect 4530 -64020 26670 -63920
<< via2 >>
rect -1070 8100 -990 8180
rect -830 8100 -750 8180
rect 3060 8110 3140 8190
rect 3280 8110 3360 8190
rect 11080 8110 11160 8190
rect 11310 8110 11390 8190
rect 15900 8100 15980 8180
rect 16140 8100 16220 8180
rect 14830 4470 14930 4570
rect 14830 4270 14930 4370
rect -1430 880 -1350 960
rect -1220 880 -1140 960
rect -1430 740 -1350 820
rect -1220 740 -1140 820
rect -270 870 -190 950
rect -50 870 30 950
rect -270 730 -190 810
rect -50 730 30 810
rect 930 900 1010 980
rect 1170 900 1250 980
rect 930 740 1010 820
rect 1170 740 1250 820
rect 18650 -2080 18730 -2000
rect 18650 -2240 18730 -2160
rect 2380 -3420 2460 -3340
rect 2540 -3420 2620 -3340
rect -2290 -4300 -2210 -4220
rect -2040 -4300 -1960 -4220
rect -2290 -4450 -2210 -4370
rect -2040 -4450 -1960 -4370
rect 13300 -3650 13380 -3570
rect 13300 -3890 13380 -3810
rect -1430 -5710 -1350 -5630
rect -1230 -5710 -1150 -5630
rect -1430 -5850 -1350 -5770
rect -1230 -5850 -1150 -5770
rect -40 -5710 40 -5630
rect 160 -5710 240 -5630
rect -40 -5850 40 -5770
rect 160 -5850 240 -5770
rect -1930 -7290 -1850 -7210
rect -1770 -7290 -1690 -7210
rect -1610 -7290 -1530 -7210
rect -1610 -9340 -1530 -9260
rect -1380 -9340 -1300 -9260
rect 610 -9340 690 -9260
rect 840 -9340 920 -9260
rect 8040 -9770 8120 -9690
rect 8260 -9770 8340 -9690
rect 18650 -7150 18730 -7070
rect 18650 -7310 18730 -7230
rect 12270 -8310 12350 -8230
rect 12510 -8310 12590 -8230
rect 16100 -9770 16180 -9690
rect 16340 -9770 16420 -9690
rect 25420 -10850 25620 -10650
rect 25820 -10850 26020 -10650
rect 26220 -10850 26420 -10650
rect 25350 -63920 25550 -63720
rect 25750 -63920 25950 -63720
rect 26150 -63920 26350 -63720
<< metal3 >>
rect -6324 11740 22100 11900
rect -6324 11640 -6240 11740
rect -6140 11640 -6040 11740
rect -5940 11730 15920 11740
rect -5940 11640 -1070 11730
rect -6324 11630 -1070 11640
rect -970 11630 -870 11730
rect -770 11630 3060 11730
rect 3160 11630 3260 11730
rect 3360 11630 11080 11730
rect 11180 11630 11280 11730
rect 11380 11640 15920 11730
rect 16020 11640 16120 11740
rect 16220 11730 22100 11740
rect 16220 11640 21620 11730
rect 11380 11630 21620 11640
rect 21720 11630 21820 11730
rect 21920 11630 22100 11730
rect -6324 11540 22100 11630
rect -6324 11440 -6240 11540
rect -6140 11440 -6040 11540
rect -5940 11530 15920 11540
rect -5940 11440 -1070 11530
rect -6324 11430 -1070 11440
rect -970 11430 -870 11530
rect -770 11430 3060 11530
rect 3160 11430 3260 11530
rect 3360 11430 11080 11530
rect 11180 11430 11280 11530
rect 11380 11440 15920 11530
rect 16020 11440 16120 11540
rect 16220 11530 22100 11540
rect 16220 11440 21620 11530
rect 11380 11430 21620 11440
rect 21720 11430 21820 11530
rect 21920 11430 22100 11530
rect -6324 11356 22100 11430
rect -4148 9740 20060 9860
rect -4148 9640 -4070 9740
rect -3970 9640 -3870 9740
rect -3770 9730 20060 9740
rect -3770 9640 19700 9730
rect -4148 9630 19700 9640
rect 19800 9630 19900 9730
rect 20000 9630 20060 9730
rect -4148 9540 20060 9630
rect -4148 9440 -4070 9540
rect -3970 9440 -3870 9540
rect -3770 9530 20060 9540
rect -3770 9440 19700 9530
rect -4148 9430 19700 9440
rect 19800 9430 19900 9530
rect 20000 9430 20060 9530
rect -4148 9316 20060 9430
rect 3020 8350 3420 8370
rect 3020 8250 3060 8350
rect 3160 8250 3260 8350
rect 3360 8250 3420 8350
rect -1110 8200 -710 8210
rect -1110 8080 -1090 8200
rect -970 8080 -850 8200
rect -730 8080 -710 8200
rect -1110 8070 -710 8080
rect 3020 8190 3420 8250
rect 3020 8110 3060 8190
rect 3140 8110 3280 8190
rect 3360 8110 3420 8190
rect 3020 8070 3420 8110
rect 11040 8350 11440 8370
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 8190 11440 8250
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8070 11440 8110
rect 15870 8330 16270 8350
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 8180 16270 8230
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8070 16270 8100
rect 14680 4570 20050 4630
rect 14680 4470 14830 4570
rect 14930 4470 19600 4570
rect 19700 4470 19900 4570
rect 20000 4470 20050 4570
rect 14680 4370 20050 4470
rect 14680 4270 14830 4370
rect 14930 4270 19600 4370
rect 19700 4270 19900 4370
rect 20000 4270 20050 4370
rect 14680 4230 20050 4270
rect -6290 1050 1290 1110
rect -6290 950 -6250 1050
rect -6150 950 -6050 1050
rect -5950 980 1290 1050
rect -5950 960 930 980
rect -5950 950 -1430 960
rect -6290 880 -1430 950
rect -1350 880 -1220 960
rect -1140 950 930 960
rect -1140 880 -270 950
rect -6290 870 -270 880
rect -190 870 -50 950
rect 30 900 930 950
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 30 870 1290 900
rect -6290 850 1290 870
rect -6290 750 -6250 850
rect -6150 750 -6050 850
rect -5950 820 1290 850
rect -5950 750 -1430 820
rect -6290 740 -1430 750
rect -1350 740 -1220 820
rect -1140 810 930 820
rect -1140 740 -270 810
rect -6290 730 -270 740
rect -190 730 -50 810
rect 30 740 930 810
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 30 730 1290 740
rect -6290 710 1290 730
rect 18510 -2000 20050 -1950
rect 18510 -2080 18650 -2000
rect 18730 -2080 19710 -2000
rect 18510 -2100 19710 -2080
rect 19810 -2100 19910 -2000
rect 20010 -2100 20050 -2000
rect 18510 -2160 20050 -2100
rect 18510 -2240 18650 -2160
rect 18730 -2200 20050 -2160
rect 18730 -2240 19710 -2200
rect 18510 -2300 19710 -2240
rect 19810 -2300 19910 -2200
rect 20010 -2300 20050 -2200
rect 18510 -2350 20050 -2300
rect -4130 -3120 2760 -3080
rect -4130 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 2760 -3120
rect -4130 -3320 2760 -3220
rect -4130 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3340 2760 -3320
rect -3770 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect -4130 -3480 2760 -3420
rect 13160 -3570 21980 -3540
rect 13160 -3650 13300 -3570
rect 13380 -3580 21980 -3570
rect 13380 -3650 21630 -3580
rect 13160 -3680 21630 -3650
rect 21730 -3680 21830 -3580
rect 21930 -3680 21980 -3580
rect 13160 -3780 21980 -3680
rect 13160 -3810 21630 -3780
rect 13160 -3890 13300 -3810
rect 13380 -3880 21630 -3810
rect 21730 -3880 21830 -3780
rect 21930 -3880 21980 -3780
rect 13380 -3890 21980 -3880
rect 13160 -3940 21980 -3890
rect -6290 -4220 -1920 -4190
rect -6290 -4230 -2290 -4220
rect -6290 -4330 -6240 -4230
rect -6140 -4330 -6040 -4230
rect -5940 -4300 -2290 -4230
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -5940 -4330 -1920 -4300
rect -6290 -4370 -1920 -4330
rect -6290 -4430 -2290 -4370
rect -6290 -4530 -6240 -4430
rect -6140 -4530 -6040 -4430
rect -5940 -4450 -2290 -4430
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -5940 -4530 -1920 -4450
rect -6290 -4590 -1920 -4530
rect -4130 -5520 310 -5470
rect -4130 -5620 -4090 -5520
rect -3990 -5620 -3890 -5520
rect -3790 -5620 310 -5520
rect -4130 -5630 310 -5620
rect -4130 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 -40 -5630
rect 40 -5710 160 -5630
rect 240 -5710 310 -5630
rect -4130 -5720 310 -5710
rect -4130 -5820 -4090 -5720
rect -3990 -5820 -3890 -5720
rect -3790 -5770 310 -5720
rect -3790 -5820 -1430 -5770
rect -4130 -5850 -1430 -5820
rect -1350 -5850 -1230 -5770
rect -1150 -5850 -40 -5770
rect 40 -5850 160 -5770
rect 240 -5850 310 -5770
rect -4130 -5870 310 -5850
rect 18510 -6990 20050 -6940
rect -4130 -7080 -1480 -7030
rect -4130 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -1480 -7080
rect -4130 -7210 -1480 -7180
rect -4130 -7280 -1930 -7210
rect -4130 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7290 -1930 -7280
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -3790 -7320 -1480 -7290
rect 18510 -7070 19700 -6990
rect 18510 -7150 18650 -7070
rect 18730 -7090 19700 -7070
rect 19800 -7090 19900 -6990
rect 20000 -7090 20050 -6990
rect 18730 -7150 20050 -7090
rect 18510 -7190 20050 -7150
rect 18510 -7230 19700 -7190
rect 18510 -7310 18650 -7230
rect 18730 -7290 19700 -7230
rect 19800 -7290 19900 -7190
rect 20000 -7290 20050 -7190
rect 18730 -7310 20050 -7290
rect -3790 -7380 -3730 -7320
rect 18510 -7340 20050 -7310
rect -4130 -7430 -3730 -7380
rect 12250 -8230 12650 -8220
rect 12250 -8310 12270 -8230
rect 12350 -8310 12510 -8230
rect 12590 -8310 12650 -8230
rect 12250 -8330 12650 -8310
rect 12250 -8430 12280 -8330
rect 12380 -8430 12480 -8330
rect 12580 -8430 12650 -8330
rect 12250 -8440 12650 -8430
rect -1640 -9260 -1240 -9240
rect -1640 -9340 -1610 -9260
rect -1530 -9340 -1380 -9260
rect -1300 -9340 -1240 -9260
rect -1640 -9380 -1240 -9340
rect -1640 -9480 -1610 -9380
rect -1510 -9480 -1410 -9380
rect -1310 -9480 -1240 -9380
rect 580 -9260 980 -9240
rect 580 -9340 610 -9260
rect 690 -9340 840 -9260
rect 920 -9340 980 -9260
rect 580 -9370 980 -9340
rect 580 -9470 600 -9370
rect 700 -9470 800 -9370
rect 900 -9470 980 -9370
rect 580 -9480 980 -9470
rect -1640 -9500 -1240 -9480
rect 8000 -9690 8390 -9660
rect 8000 -9770 8040 -9690
rect 8120 -9770 8260 -9690
rect 8340 -9770 8390 -9690
rect 8000 -9800 8390 -9770
rect 8000 -9900 8030 -9800
rect 8130 -9900 8250 -9800
rect 8350 -9900 8390 -9800
rect 8000 -9910 8390 -9900
rect 16070 -9690 16460 -9660
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9820 16460 -9770
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -9940 16460 -9920
rect 25228 -10650 26860 -10404
rect 25228 -10850 25420 -10650
rect 25620 -10850 25820 -10650
rect 26020 -10850 26220 -10650
rect 26420 -10850 26860 -10650
rect 25228 -11084 26860 -10850
rect -4148 -11510 20060 -11356
rect -4148 -11610 -4070 -11510
rect -3970 -11610 -3870 -11510
rect -3770 -11520 20060 -11510
rect -3770 -11610 8040 -11520
rect -4148 -11620 8040 -11610
rect 8140 -11620 8240 -11520
rect 8340 -11620 16120 -11520
rect 16220 -11620 16320 -11520
rect 16420 -11530 20060 -11520
rect 16420 -11620 19690 -11530
rect -4148 -11630 19690 -11620
rect 19790 -11630 19890 -11530
rect 19990 -11630 20060 -11530
rect -4148 -11710 20060 -11630
rect -4148 -11810 -4070 -11710
rect -3970 -11810 -3870 -11710
rect -3770 -11720 20060 -11710
rect -3770 -11810 8040 -11720
rect -4148 -11820 8040 -11810
rect 8140 -11820 8240 -11720
rect 8340 -11820 16120 -11720
rect 16220 -11820 16320 -11720
rect 16420 -11730 20060 -11720
rect 16420 -11820 19690 -11730
rect -4148 -11830 19690 -11820
rect 19790 -11830 19890 -11730
rect 19990 -11830 20060 -11730
rect -4148 -11900 20060 -11830
rect -6324 -13710 22100 -13532
rect -6324 -13720 630 -13710
rect -6324 -13820 -6240 -13720
rect -6140 -13820 -6040 -13720
rect -5940 -13730 630 -13720
rect -5940 -13820 -1600 -13730
rect -6324 -13830 -1600 -13820
rect -1500 -13830 -1400 -13730
rect -1300 -13810 630 -13730
rect 730 -13810 830 -13710
rect 930 -13810 12300 -13710
rect 12400 -13810 12500 -13710
rect 12600 -13730 22100 -13710
rect 12600 -13810 21620 -13730
rect -1300 -13830 21620 -13810
rect 21720 -13830 21820 -13730
rect 21920 -13830 22100 -13730
rect -6324 -13910 22100 -13830
rect -6324 -13920 630 -13910
rect -6324 -14020 -6240 -13920
rect -6140 -14020 -6040 -13920
rect -5940 -13930 630 -13920
rect -5940 -14020 -1600 -13930
rect -6324 -14030 -1600 -14020
rect -1500 -14030 -1400 -13930
rect -1300 -14010 630 -13930
rect 730 -14010 830 -13910
rect 930 -14010 12300 -13910
rect 12400 -14010 12500 -13910
rect 12600 -13930 22100 -13910
rect 12600 -14010 21620 -13930
rect -1300 -14030 21620 -14010
rect 21720 -14030 21820 -13930
rect 21920 -14030 22100 -13930
rect -6324 -14076 22100 -14030
rect 25092 -63720 26724 -63580
rect 25092 -63920 25350 -63720
rect 25550 -63920 25750 -63720
rect 25950 -63920 26150 -63720
rect 26350 -63920 26724 -63720
rect 25092 -64124 26724 -63920
<< via3 >>
rect -6240 11640 -6140 11740
rect -6040 11640 -5940 11740
rect -1070 11630 -970 11730
rect -870 11630 -770 11730
rect 3060 11630 3160 11730
rect 3260 11630 3360 11730
rect 11080 11630 11180 11730
rect 11280 11630 11380 11730
rect 15920 11640 16020 11740
rect 16120 11640 16220 11740
rect 21620 11630 21720 11730
rect 21820 11630 21920 11730
rect -6240 11440 -6140 11540
rect -6040 11440 -5940 11540
rect -1070 11430 -970 11530
rect -870 11430 -770 11530
rect 3060 11430 3160 11530
rect 3260 11430 3360 11530
rect 11080 11430 11180 11530
rect 11280 11430 11380 11530
rect 15920 11440 16020 11540
rect 16120 11440 16220 11540
rect 21620 11430 21720 11530
rect 21820 11430 21920 11530
rect -4070 9640 -3970 9740
rect -3870 9640 -3770 9740
rect 19700 9630 19800 9730
rect 19900 9630 20000 9730
rect -4070 9440 -3970 9540
rect -3870 9440 -3770 9540
rect 19700 9430 19800 9530
rect 19900 9430 20000 9530
rect 3060 8250 3160 8350
rect 3260 8250 3360 8350
rect -1090 8180 -970 8200
rect -1090 8100 -1070 8180
rect -1070 8100 -990 8180
rect -990 8100 -970 8180
rect -1090 8080 -970 8100
rect -850 8180 -730 8200
rect -850 8100 -830 8180
rect -830 8100 -750 8180
rect -750 8100 -730 8180
rect -850 8080 -730 8100
rect 11080 8250 11180 8350
rect 11280 8250 11380 8350
rect 15900 8230 16000 8330
rect 16130 8230 16230 8330
rect 19600 4470 19700 4570
rect 19900 4470 20000 4570
rect 19600 4270 19700 4370
rect 19900 4270 20000 4370
rect -6250 950 -6150 1050
rect -6050 950 -5950 1050
rect -6250 750 -6150 850
rect -6050 750 -5950 850
rect 19710 -2100 19810 -2000
rect 19910 -2100 20010 -2000
rect 19710 -2300 19810 -2200
rect 19910 -2300 20010 -2200
rect -4070 -3220 -3970 -3120
rect -3870 -3220 -3770 -3120
rect -4070 -3420 -3970 -3320
rect -3870 -3420 -3770 -3320
rect 21630 -3680 21730 -3580
rect 21830 -3680 21930 -3580
rect 21630 -3880 21730 -3780
rect 21830 -3880 21930 -3780
rect -6240 -4330 -6140 -4230
rect -6040 -4330 -5940 -4230
rect -6240 -4530 -6140 -4430
rect -6040 -4530 -5940 -4430
rect -4090 -5620 -3990 -5520
rect -3890 -5620 -3790 -5520
rect -4090 -5820 -3990 -5720
rect -3890 -5820 -3790 -5720
rect -4090 -7180 -3990 -7080
rect -3890 -7180 -3790 -7080
rect -4090 -7380 -3990 -7280
rect -3890 -7380 -3790 -7280
rect 19700 -7090 19800 -6990
rect 19900 -7090 20000 -6990
rect 19700 -7290 19800 -7190
rect 19900 -7290 20000 -7190
rect 12280 -8430 12380 -8330
rect 12480 -8430 12580 -8330
rect -1610 -9480 -1510 -9380
rect -1410 -9480 -1310 -9380
rect 600 -9470 700 -9370
rect 800 -9470 900 -9370
rect 8030 -9900 8130 -9800
rect 8250 -9900 8350 -9800
rect 16110 -9920 16210 -9820
rect 16310 -9920 16410 -9820
rect -4070 -11610 -3970 -11510
rect -3870 -11610 -3770 -11510
rect 8040 -11620 8140 -11520
rect 8240 -11620 8340 -11520
rect 16120 -11620 16220 -11520
rect 16320 -11620 16420 -11520
rect 19690 -11630 19790 -11530
rect 19890 -11630 19990 -11530
rect -4070 -11810 -3970 -11710
rect -3870 -11810 -3770 -11710
rect 8040 -11820 8140 -11720
rect 8240 -11820 8340 -11720
rect 16120 -11820 16220 -11720
rect 16320 -11820 16420 -11720
rect 19690 -11830 19790 -11730
rect 19890 -11830 19990 -11730
rect -6240 -13820 -6140 -13720
rect -6040 -13820 -5940 -13720
rect -1600 -13830 -1500 -13730
rect -1400 -13830 -1300 -13730
rect 630 -13810 730 -13710
rect 830 -13810 930 -13710
rect 12300 -13810 12400 -13710
rect 12500 -13810 12600 -13710
rect 21620 -13830 21720 -13730
rect 21820 -13830 21920 -13730
rect -6240 -14020 -6140 -13920
rect -6040 -14020 -5940 -13920
rect -1600 -14030 -1500 -13930
rect -1400 -14030 -1300 -13930
rect 630 -14010 730 -13910
rect 830 -14010 930 -13910
rect 12300 -14010 12400 -13910
rect 12500 -14010 12600 -13910
rect 21620 -14030 21720 -13930
rect 21820 -14030 21920 -13930
<< metal4 >>
rect -6324 11740 -5780 11900
rect -6324 11640 -6240 11740
rect -6140 11640 -6040 11740
rect -5940 11640 -5780 11740
rect -6324 11540 -5780 11640
rect -6324 11440 -6240 11540
rect -6140 11440 -6040 11540
rect -5940 11440 -5780 11540
rect -6324 1050 -5780 11440
rect -1110 11730 -710 11790
rect -1110 11630 -1070 11730
rect -970 11630 -870 11730
rect -770 11630 -710 11730
rect -1110 11530 -710 11630
rect -1110 11430 -1070 11530
rect -970 11430 -870 11530
rect -770 11430 -710 11530
rect -6324 950 -6250 1050
rect -6150 950 -6050 1050
rect -5950 950 -5780 1050
rect -6324 850 -5780 950
rect -6324 750 -6250 850
rect -6150 750 -6050 850
rect -5950 750 -5780 850
rect -6324 -4230 -5780 750
rect -6324 -4330 -6240 -4230
rect -6140 -4330 -6040 -4230
rect -5940 -4330 -5780 -4230
rect -6324 -4430 -5780 -4330
rect -6324 -4530 -6240 -4430
rect -6140 -4530 -6040 -4430
rect -5940 -4530 -5780 -4430
rect -6324 -13720 -5780 -4530
rect -4148 9740 -3604 9860
rect -4148 9640 -4070 9740
rect -3970 9640 -3870 9740
rect -3770 9640 -3604 9740
rect -4148 9540 -3604 9640
rect -4148 9440 -4070 9540
rect -3970 9440 -3870 9540
rect -3770 9440 -3604 9540
rect -4148 -3120 -3604 9440
rect -1110 8200 -710 11430
rect -1110 8080 -1090 8200
rect -970 8080 -850 8200
rect -730 8080 -710 8200
rect -1110 7990 -710 8080
rect 3020 11730 3420 11790
rect 3020 11630 3060 11730
rect 3160 11630 3260 11730
rect 3360 11630 3420 11730
rect 3020 11530 3420 11630
rect 3020 11430 3060 11530
rect 3160 11430 3260 11530
rect 3360 11430 3420 11530
rect 3020 8350 3420 11430
rect 3020 8250 3060 8350
rect 3160 8250 3260 8350
rect 3360 8250 3420 8350
rect 3020 7990 3420 8250
rect 11040 11730 11440 11790
rect 11040 11630 11080 11730
rect 11180 11630 11280 11730
rect 11380 11630 11440 11730
rect 11040 11530 11440 11630
rect 11040 11430 11080 11530
rect 11180 11430 11280 11530
rect 11380 11430 11440 11530
rect 11040 8350 11440 11430
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 7990 11440 8250
rect 15870 11740 16270 11790
rect 15870 11640 15920 11740
rect 16020 11640 16120 11740
rect 16220 11640 16270 11740
rect 15870 11540 16270 11640
rect 15870 11440 15920 11540
rect 16020 11440 16120 11540
rect 16220 11440 16270 11540
rect 15870 8330 16270 11440
rect 21556 11730 22100 11900
rect 21556 11630 21620 11730
rect 21720 11630 21820 11730
rect 21920 11630 22100 11730
rect 21556 11530 22100 11630
rect 21556 11430 21620 11530
rect 21720 11430 21820 11530
rect 21920 11430 22100 11530
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 7990 16270 8230
rect 19516 9730 20060 9860
rect 19516 9630 19700 9730
rect 19800 9630 19900 9730
rect 20000 9630 20060 9730
rect 19516 9530 20060 9630
rect 19516 9430 19700 9530
rect 19800 9430 19900 9530
rect 20000 9430 20060 9530
rect -4148 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 -3604 -3120
rect -4148 -3320 -3604 -3220
rect -4148 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3420 -3604 -3320
rect -4148 -5520 -3604 -3420
rect -4148 -5620 -4090 -5520
rect -3990 -5620 -3890 -5520
rect -3790 -5620 -3604 -5520
rect -4148 -5720 -3604 -5620
rect -4148 -5820 -4090 -5720
rect -3990 -5820 -3890 -5720
rect -3790 -5820 -3604 -5720
rect -4148 -7080 -3604 -5820
rect -4148 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -3604 -7080
rect -4148 -7280 -3604 -7180
rect -4148 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7380 -3604 -7280
rect -4148 -11510 -3604 -7380
rect 19516 4570 20060 9430
rect 19516 4470 19600 4570
rect 19700 4470 19900 4570
rect 20000 4470 20060 4570
rect 19516 4370 20060 4470
rect 19516 4270 19600 4370
rect 19700 4270 19900 4370
rect 20000 4270 20060 4370
rect 19516 -2000 20060 4270
rect 19516 -2100 19710 -2000
rect 19810 -2100 19910 -2000
rect 20010 -2100 20060 -2000
rect 19516 -2200 20060 -2100
rect 19516 -2300 19710 -2200
rect 19810 -2300 19910 -2200
rect 20010 -2300 20060 -2200
rect 19516 -6990 20060 -2300
rect 19516 -7090 19700 -6990
rect 19800 -7090 19900 -6990
rect 20000 -7090 20060 -6990
rect 19516 -7190 20060 -7090
rect 19516 -7290 19700 -7190
rect 19800 -7290 19900 -7190
rect 20000 -7290 20060 -7190
rect 12250 -8330 12650 -8120
rect 12250 -8430 12280 -8330
rect 12380 -8430 12480 -8330
rect 12580 -8430 12650 -8330
rect -4148 -11610 -4070 -11510
rect -3970 -11610 -3870 -11510
rect -3770 -11610 -3604 -11510
rect -4148 -11710 -3604 -11610
rect -4148 -11810 -4070 -11710
rect -3970 -11810 -3870 -11710
rect -3770 -11810 -3604 -11710
rect -4148 -11900 -3604 -11810
rect -1640 -9380 -1240 -9150
rect -1640 -9480 -1610 -9380
rect -1510 -9480 -1410 -9380
rect -1310 -9480 -1240 -9380
rect -6324 -13820 -6240 -13720
rect -6140 -13820 -6040 -13720
rect -5940 -13820 -5780 -13720
rect -6324 -13920 -5780 -13820
rect -6324 -14020 -6240 -13920
rect -6140 -14020 -6040 -13920
rect -5940 -14020 -5780 -13920
rect -6324 -14076 -5780 -14020
rect -1640 -13730 -1240 -9480
rect -1640 -13830 -1600 -13730
rect -1500 -13830 -1400 -13730
rect -1300 -13830 -1240 -13730
rect -1640 -13930 -1240 -13830
rect -1640 -14030 -1600 -13930
rect -1500 -14030 -1400 -13930
rect -1300 -14030 -1240 -13930
rect -1640 -14070 -1240 -14030
rect 580 -9370 980 -9140
rect 580 -9470 600 -9370
rect 700 -9470 800 -9370
rect 900 -9470 980 -9370
rect 580 -13710 980 -9470
rect 8000 -9800 8390 -9550
rect 8000 -9900 8030 -9800
rect 8130 -9900 8250 -9800
rect 8350 -9900 8390 -9800
rect 8000 -11520 8390 -9900
rect 8000 -11620 8040 -11520
rect 8140 -11620 8240 -11520
rect 8340 -11620 8390 -11520
rect 8000 -11720 8390 -11620
rect 8000 -11820 8040 -11720
rect 8140 -11820 8240 -11720
rect 8340 -11820 8390 -11720
rect 8000 -11870 8390 -11820
rect 580 -13810 630 -13710
rect 730 -13810 830 -13710
rect 930 -13810 980 -13710
rect 580 -13910 980 -13810
rect 580 -14010 630 -13910
rect 730 -14010 830 -13910
rect 930 -14010 980 -13910
rect 580 -14070 980 -14010
rect 12250 -13710 12650 -8430
rect 16070 -9820 16460 -9560
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -11520 16460 -9920
rect 16070 -11620 16120 -11520
rect 16220 -11620 16320 -11520
rect 16420 -11620 16460 -11520
rect 16070 -11720 16460 -11620
rect 16070 -11820 16120 -11720
rect 16220 -11820 16320 -11720
rect 16420 -11820 16460 -11720
rect 16070 -11870 16460 -11820
rect 19516 -11530 20060 -7290
rect 19516 -11630 19690 -11530
rect 19790 -11630 19890 -11530
rect 19990 -11630 20060 -11530
rect 19516 -11730 20060 -11630
rect 19516 -11830 19690 -11730
rect 19790 -11830 19890 -11730
rect 19990 -11830 20060 -11730
rect 19516 -11900 20060 -11830
rect 21556 -3580 22100 11430
rect 21556 -3680 21630 -3580
rect 21730 -3680 21830 -3580
rect 21930 -3680 22100 -3580
rect 21556 -3780 22100 -3680
rect 21556 -3880 21630 -3780
rect 21730 -3880 21830 -3780
rect 21930 -3880 22100 -3780
rect 12250 -13810 12300 -13710
rect 12400 -13810 12500 -13710
rect 12600 -13810 12650 -13710
rect 12250 -13910 12650 -13810
rect 12250 -14010 12300 -13910
rect 12400 -14010 12500 -13910
rect 12600 -14010 12650 -13910
rect 12250 -14070 12650 -14010
rect 21556 -13730 22100 -3880
rect 21556 -13830 21620 -13730
rect 21720 -13830 21820 -13730
rect 21920 -13830 22100 -13730
rect 21556 -13930 22100 -13830
rect 21556 -14030 21620 -13930
rect 21720 -14030 21820 -13930
rect 21920 -14030 22100 -13930
rect 21556 -14076 22100 -14030
use ALib_DCO  ALib_DCO_0 ./../dco
timestamp 1730531556
transform 1 0 5200 0 1 -5190
box 1000 -4470 13410 5980
use ALib_VCO  ALib_VCO_0 ./../vco
timestamp 1730639796
transform 1 0 -2020 0 1 1040
box 0 280 20640 7030
use DLib_Quantizer  DLib_Quantizer_0 ./../quantizer
timestamp 1730532965
transform 1 0 -2210 0 1 -4630
box 190 -710 5890 730
use DLib_UpDownCounter  DLib_UpDownCounter_0 ./../count
timestamp 1730536752
transform 1 0 -1140 0 1 -5986
box -880 -3154 3140 -440
use DLib_UpDownCounter  DLib_UpDownCounter_1
timestamp 1730536752
transform 1 0 -1140 0 1 344
box -880 -3154 3140 -440
<< labels >>
flabel metal3 -5940 11356 -1070 11900 1 FreeSans 2176 0 0 0 VDDA
port 7 nsew power input
flabel metal3 16388 9316 19516 9860 1 FreeSans 2176 0 0 0 GND
port 8 nsew ground input
flabel metal3 25092 -64124 26724 -63580 1 FreeSans 1088 0 0 0 Vbs_12
port 1 nsew signal input
flabel metal3 25228 -11084 26860 -10404 1 FreeSans 1088 0 0 0 Vbs_34
port 2 nsew signal input
flabel metal2 17342 34914 17710 36938 1 FreeSans 736 0 0 0 Anlg_in
port 3 nsew signal input
flabel metal2 -7590 -17526 -7038 -16330 1 FreeSans 736 0 0 0 ENB
port 4 nsew signal input
flabel metal2 -5198 -17526 -4646 -16330 1 FreeSans 736 0 0 0 CLK
port 5 nsew signal input
flabel metal2 2806 -17526 3358 -16330 1 FreeSans 736 0 0 0 Dout
port 6 nsew signal input
<< end >>
