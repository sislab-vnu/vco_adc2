magic
tech sky130A
timestamp 1730541949
<< locali >>
rect 565 -780 3055 -770
rect 565 -800 575 -780
rect 595 -800 615 -780
rect 635 -800 2985 -780
rect 3005 -800 3025 -780
rect 3045 -800 3055 -780
rect 565 -810 3055 -800
rect 3015 -820 3055 -810
rect 3015 -840 3025 -820
rect 3045 -840 3055 -820
rect 3015 -850 3055 -840
rect 735 -1075 1370 -1065
rect 735 -1105 1210 -1075
rect 1240 -1105 1270 -1075
rect 1300 -1105 1330 -1075
rect 1360 -1105 1370 -1075
rect 735 -1110 1370 -1105
rect 765 -1115 1370 -1110
rect -1120 -3375 -915 -3370
rect -1120 -3380 -910 -3375
rect -1120 -3400 -1110 -3380
rect -1090 -3400 -1070 -3380
rect -1050 -3400 -910 -3380
rect -1120 -3410 -910 -3400
rect -1120 -3420 -1080 -3410
rect -1120 -3440 -1110 -3420
rect -1090 -3440 -1080 -3420
rect -1120 -3450 -1080 -3440
rect 630 -3945 1185 -3935
rect 630 -3965 640 -3945
rect 660 -3965 680 -3945
rect 700 -3965 720 -3945
rect 740 -3965 1075 -3945
rect 1095 -3965 1115 -3945
rect 1135 -3965 1155 -3945
rect 1175 -3965 1185 -3945
rect 630 -3975 1185 -3965
rect 8140 -3950 8585 -3935
rect 8140 -3970 8155 -3950
rect 8175 -3970 8195 -3950
rect 8215 -3970 8585 -3950
rect 8140 -3985 8585 -3970
rect 8140 -3990 8190 -3985
rect 8140 -4010 8155 -3990
rect 8175 -4010 8190 -3990
rect 8140 -4025 8190 -4010
rect 8535 -4980 8585 -3985
rect 8535 -5000 8550 -4980
rect 8570 -5000 8585 -4980
rect 8535 -5010 8585 -5000
rect 8500 -5020 8585 -5010
rect 8500 -5040 8510 -5020
rect 8530 -5040 8550 -5020
rect 8570 -5040 8585 -5020
rect 8500 -5050 8585 -5040
<< viali >>
rect -545 4005 -525 4025
rect -505 4005 -485 4025
rect -465 4005 -445 4025
rect -425 4005 -405 4025
rect -385 4005 -365 4025
rect 1520 4005 1540 4025
rect 1560 4005 1580 4025
rect 1600 4005 1620 4025
rect 1640 4005 1660 4025
rect 1680 4005 1700 4025
rect 5530 4005 5550 4025
rect 5570 4005 5590 4025
rect 5610 4005 5630 4025
rect 5650 4005 5670 4025
rect 5690 4005 5710 4025
rect 7945 4005 7965 4025
rect 7985 4005 8005 4025
rect 8025 4005 8045 4025
rect 8065 4005 8085 4025
rect 8105 4005 8125 4025
rect -1000 -235 -980 -215
rect -960 -235 -940 -215
rect 575 -800 595 -780
rect 615 -800 635 -780
rect 2985 -800 3005 -780
rect 3025 -800 3045 -780
rect 3025 -840 3045 -820
rect 1210 -1105 1240 -1075
rect 1270 -1105 1300 -1075
rect 1330 -1105 1360 -1075
rect -1110 -3400 -1090 -3380
rect -1070 -3400 -1050 -3380
rect -1110 -3440 -1090 -3420
rect 640 -3965 660 -3945
rect 680 -3965 700 -3945
rect 720 -3965 740 -3945
rect 1075 -3965 1095 -3945
rect 1115 -3965 1135 -3945
rect 1155 -3965 1175 -3945
rect 8155 -3970 8175 -3950
rect 8195 -3970 8215 -3950
rect 8155 -4010 8175 -3990
rect 8550 -5000 8570 -4980
rect 8510 -5040 8530 -5020
rect 8550 -5040 8570 -5020
<< metal1 >>
rect -555 4030 -355 4035
rect -555 4000 -550 4030
rect -520 4025 -490 4030
rect -460 4025 -430 4030
rect -400 4025 -355 4030
rect -520 4005 -505 4025
rect -445 4005 -430 4025
rect -400 4005 -385 4025
rect -365 4005 -355 4025
rect -520 4000 -490 4005
rect -460 4000 -430 4005
rect -400 4000 -355 4005
rect -555 3995 -355 4000
rect 1510 4030 1710 4035
rect 1510 4000 1515 4030
rect 1545 4025 1595 4030
rect 1625 4025 1675 4030
rect 1545 4005 1560 4025
rect 1580 4005 1595 4025
rect 1625 4005 1640 4025
rect 1660 4005 1675 4025
rect 1545 4000 1595 4005
rect 1625 4000 1675 4005
rect 1705 4000 1710 4030
rect 1510 3995 1710 4000
rect 5520 4030 5720 4035
rect 5520 4000 5525 4030
rect 5555 4025 5605 4030
rect 5635 4025 5685 4030
rect 5555 4005 5570 4025
rect 5590 4005 5605 4025
rect 5635 4005 5650 4025
rect 5670 4005 5685 4025
rect 5555 4000 5605 4005
rect 5635 4000 5685 4005
rect 5715 4000 5720 4030
rect 5520 3995 5720 4000
rect 7935 4030 8135 4035
rect 7935 4000 7940 4030
rect 7970 4025 8020 4030
rect 8050 4025 8100 4030
rect 7970 4005 7985 4025
rect 8005 4005 8020 4025
rect 8050 4005 8065 4025
rect 8085 4005 8100 4025
rect 7970 4000 8020 4005
rect 8050 4000 8100 4005
rect 8130 4000 8135 4030
rect 7935 3995 8135 4000
rect -1010 -205 -960 1050
rect -740 540 -540 555
rect -740 505 -715 540
rect -680 505 -600 540
rect -565 505 -540 540
rect -740 -65 -540 505
rect -160 535 40 555
rect -160 500 -135 535
rect -100 500 -25 535
rect 10 500 40 535
rect -160 -60 40 500
rect 445 540 645 555
rect 445 510 465 540
rect 495 510 590 540
rect 620 510 645 540
rect 445 -65 645 510
rect -1010 -215 -930 -205
rect -1010 -235 -1000 -215
rect -980 -235 -960 -215
rect -940 -235 -930 -215
rect -1010 -245 -930 -235
rect 485 -780 645 -770
rect 485 -800 575 -780
rect 595 -800 615 -780
rect 635 -800 645 -780
rect 485 -810 645 -800
rect 2975 -780 3055 -770
rect 2975 -800 2985 -780
rect 3005 -800 3025 -780
rect 3045 -800 3055 -780
rect 2975 -810 3055 -800
rect 3015 -820 3055 -810
rect 3015 -840 3025 -820
rect 3045 -840 3055 -820
rect 1200 -1075 1370 -1065
rect 1200 -1105 1210 -1075
rect 1240 -1105 1270 -1075
rect 1300 -1105 1330 -1075
rect 1360 -1105 1370 -1075
rect 1200 -1115 1370 -1105
rect 1180 -1550 1380 -1115
rect 1180 -1580 1195 -1550
rect 1225 -1580 1255 -1550
rect 1285 -1580 1315 -1550
rect 1345 -1580 1380 -1550
rect 1180 -1610 1380 -1580
rect 1180 -1640 1195 -1610
rect 1225 -1640 1255 -1610
rect 1285 -1640 1315 -1610
rect 1345 -1640 1380 -1610
rect 1180 -1740 1380 -1640
rect -1160 -2245 -960 -1950
rect -1160 -2275 -1140 -2245
rect -1110 -2275 -1015 -2245
rect -985 -2275 -960 -2245
rect -1160 -2400 -960 -2275
rect 3015 -2415 3055 -840
rect 6580 -1790 6625 -1770
rect 6580 -1820 6585 -1790
rect 6615 -1820 6625 -1790
rect 6580 -1850 6625 -1820
rect 6580 -1880 6585 -1850
rect 6615 -1880 6625 -1850
rect 6580 -1945 6625 -1880
rect 3015 -2455 3260 -2415
rect -895 -3035 -855 -2510
rect -740 -2750 -540 -2670
rect -740 -2780 -725 -2750
rect -695 -2780 -665 -2750
rect -635 -2780 -605 -2750
rect -575 -2780 -540 -2750
rect -740 -2790 -540 -2780
rect -895 -3075 1185 -3035
rect -1120 -3380 -1040 -3370
rect -1120 -3400 -1110 -3380
rect -1090 -3400 -1070 -3380
rect -1050 -3400 -1040 -3380
rect -1120 -3410 -1040 -3400
rect -1120 -3420 -1080 -3410
rect -1120 -3440 -1110 -3420
rect -1090 -3440 -1080 -3420
rect -1120 -5010 -1080 -3440
rect -980 -3545 -740 -3530
rect -980 -3575 -965 -3545
rect -935 -3575 -905 -3545
rect -875 -3575 -845 -3545
rect -815 -3575 -785 -3545
rect -755 -3575 -740 -3545
rect -980 -3585 -740 -3575
rect 1145 -3935 1185 -3075
rect 3220 -3505 3260 -2455
rect 485 -3945 750 -3935
rect 485 -3965 640 -3945
rect 660 -3965 680 -3945
rect 700 -3965 720 -3945
rect 740 -3965 750 -3945
rect 485 -3975 750 -3965
rect 1065 -3945 1185 -3935
rect 1065 -3965 1075 -3945
rect 1095 -3965 1115 -3945
rect 1135 -3965 1155 -3945
rect 1175 -3965 1185 -3945
rect 1065 -3975 1185 -3965
rect 8140 -3950 8245 -3935
rect 8140 -3970 8155 -3950
rect 8175 -3970 8195 -3950
rect 8215 -3970 8245 -3950
rect 8140 -3985 8245 -3970
rect 8140 -3990 8190 -3985
rect 8140 -4010 8155 -3990
rect 8175 -4010 8190 -3990
rect 8140 -4025 8190 -4010
rect 6125 -4070 6325 -4060
rect 6125 -4100 6140 -4070
rect 6170 -4100 6200 -4070
rect 6230 -4100 6260 -4070
rect 6290 -4100 6325 -4070
rect 6125 -4110 6325 -4100
rect -820 -4585 -620 -4525
rect -820 -4615 -805 -4585
rect -775 -4615 -745 -4585
rect -715 -4615 -685 -4585
rect -655 -4615 -620 -4585
rect -820 -4685 -620 -4615
rect 290 -4580 490 -4530
rect 290 -4610 305 -4580
rect 335 -4610 365 -4580
rect 395 -4610 425 -4580
rect 455 -4610 490 -4580
rect 290 -4625 490 -4610
rect 8535 -4980 8585 -4970
rect 8535 -5000 8550 -4980
rect 8570 -5000 8585 -4980
rect 8535 -5010 8585 -5000
rect -1120 -5020 8585 -5010
rect -1120 -5040 8510 -5020
rect 8530 -5040 8550 -5020
rect 8570 -5040 8585 -5020
rect -1120 -5050 8585 -5040
<< via1 >>
rect -550 4025 -520 4030
rect -490 4025 -460 4030
rect -430 4025 -400 4030
rect -550 4005 -545 4025
rect -545 4005 -525 4025
rect -525 4005 -520 4025
rect -490 4005 -485 4025
rect -485 4005 -465 4025
rect -465 4005 -460 4025
rect -430 4005 -425 4025
rect -425 4005 -405 4025
rect -405 4005 -400 4025
rect -550 4000 -520 4005
rect -490 4000 -460 4005
rect -430 4000 -400 4005
rect 1515 4025 1545 4030
rect 1595 4025 1625 4030
rect 1675 4025 1705 4030
rect 1515 4005 1520 4025
rect 1520 4005 1540 4025
rect 1540 4005 1545 4025
rect 1595 4005 1600 4025
rect 1600 4005 1620 4025
rect 1620 4005 1625 4025
rect 1675 4005 1680 4025
rect 1680 4005 1700 4025
rect 1700 4005 1705 4025
rect 1515 4000 1545 4005
rect 1595 4000 1625 4005
rect 1675 4000 1705 4005
rect 5525 4025 5555 4030
rect 5605 4025 5635 4030
rect 5685 4025 5715 4030
rect 5525 4005 5530 4025
rect 5530 4005 5550 4025
rect 5550 4005 5555 4025
rect 5605 4005 5610 4025
rect 5610 4005 5630 4025
rect 5630 4005 5635 4025
rect 5685 4005 5690 4025
rect 5690 4005 5710 4025
rect 5710 4005 5715 4025
rect 5525 4000 5555 4005
rect 5605 4000 5635 4005
rect 5685 4000 5715 4005
rect 7940 4025 7970 4030
rect 8020 4025 8050 4030
rect 8100 4025 8130 4030
rect 7940 4005 7945 4025
rect 7945 4005 7965 4025
rect 7965 4005 7970 4025
rect 8020 4005 8025 4025
rect 8025 4005 8045 4025
rect 8045 4005 8050 4025
rect 8100 4005 8105 4025
rect 8105 4005 8125 4025
rect 8125 4005 8130 4025
rect 7940 4000 7970 4005
rect 8020 4000 8050 4005
rect 8100 4000 8130 4005
rect 7350 2370 7380 2400
rect 7350 2310 7380 2340
rect 7350 2250 7380 2280
rect -715 505 -680 540
rect -600 505 -565 540
rect -135 500 -100 535
rect -25 500 10 535
rect 465 510 495 540
rect 590 510 620 540
rect 1195 -1580 1225 -1550
rect 1255 -1580 1285 -1550
rect 1315 -1580 1345 -1550
rect 1195 -1640 1225 -1610
rect 1255 -1640 1285 -1610
rect 1315 -1640 1345 -1610
rect -1140 -2275 -1110 -2245
rect -1015 -2275 -985 -2245
rect 9265 -1040 9295 -1010
rect 9265 -1100 9295 -1070
rect 9265 -1160 9295 -1130
rect 6585 -1820 6615 -1790
rect 6585 -1880 6615 -1850
rect -725 -2780 -695 -2750
rect -665 -2780 -635 -2750
rect -605 -2780 -575 -2750
rect -965 -3575 -935 -3545
rect -905 -3575 -875 -3545
rect -845 -3575 -815 -3545
rect -785 -3575 -755 -3545
rect 9265 -3535 9295 -3505
rect 9265 -3595 9295 -3565
rect 9265 -3655 9295 -3625
rect 6140 -4100 6170 -4070
rect 6200 -4100 6230 -4070
rect 6260 -4100 6290 -4070
rect -805 -4615 -775 -4585
rect -745 -4615 -715 -4585
rect -685 -4615 -655 -4585
rect 305 -4610 335 -4580
rect 365 -4610 395 -4580
rect 425 -4610 455 -4580
rect 4015 -4820 4045 -4790
rect 4075 -4820 4105 -4790
rect 4135 -4820 4165 -4790
rect 8045 -4820 8075 -4790
rect 8105 -4820 8135 -4790
rect 8165 -4820 8195 -4790
<< metal2 >>
rect -555 4090 -355 4105
rect -555 4050 -535 4090
rect -495 4050 -415 4090
rect -375 4050 -355 4090
rect -555 4030 -355 4050
rect -555 4000 -550 4030
rect -520 4000 -490 4030
rect -460 4000 -430 4030
rect -400 4000 -355 4030
rect -555 3995 -355 4000
rect 1510 4095 1710 4105
rect 1510 4055 1530 4095
rect 1570 4055 1640 4095
rect 1680 4055 1710 4095
rect 1510 4030 1710 4055
rect 1510 4000 1515 4030
rect 1545 4000 1595 4030
rect 1625 4000 1675 4030
rect 1705 4000 1710 4030
rect 1510 3995 1710 4000
rect 5520 4095 5720 4110
rect 5520 4055 5540 4095
rect 5580 4055 5655 4095
rect 5695 4055 5720 4095
rect 5520 4030 5720 4055
rect 5520 4000 5525 4030
rect 5555 4000 5605 4030
rect 5635 4000 5685 4030
rect 5715 4000 5720 4030
rect 5520 3995 5720 4000
rect 7935 4090 8135 4105
rect 7935 4050 7950 4090
rect 7990 4050 8070 4090
rect 8110 4050 8135 4090
rect 7935 4030 8135 4050
rect 7935 4000 7940 4030
rect 7970 4000 8020 4030
rect 8050 4000 8100 4030
rect 8130 4000 8135 4030
rect 7935 3995 8135 4000
rect 7340 2405 7495 2435
rect 7340 2400 7415 2405
rect 7340 2370 7350 2400
rect 7380 2370 7415 2400
rect 7340 2355 7415 2370
rect 7465 2355 7495 2405
rect 7340 2340 7495 2355
rect 7340 2310 7350 2340
rect 7380 2310 7495 2340
rect 7340 2305 7495 2310
rect 7340 2280 7415 2305
rect 7340 2250 7350 2280
rect 7380 2255 7415 2280
rect 7465 2255 7495 2305
rect 7380 2250 7495 2255
rect 7340 2235 7495 2250
rect -740 540 -540 555
rect -740 505 -715 540
rect -680 505 -600 540
rect -565 505 -540 540
rect -740 480 -540 505
rect -740 440 -715 480
rect -675 440 -610 480
rect -570 440 -540 480
rect -740 410 -540 440
rect -740 370 -715 410
rect -675 370 -610 410
rect -570 370 -540 410
rect -740 355 -540 370
rect -160 535 40 555
rect -160 500 -135 535
rect -100 500 -25 535
rect 10 500 40 535
rect -160 475 40 500
rect -160 435 -135 475
rect -95 435 -25 475
rect 15 435 40 475
rect -160 405 40 435
rect -160 365 -135 405
rect -95 365 -25 405
rect 15 365 40 405
rect -160 355 40 365
rect 445 540 645 555
rect 445 510 465 540
rect 495 510 590 540
rect 620 510 645 540
rect 445 490 645 510
rect 445 450 465 490
rect 505 450 585 490
rect 625 450 645 490
rect 445 410 645 450
rect 445 370 465 410
rect 505 370 585 410
rect 625 370 645 410
rect 445 355 645 370
rect 9255 -1000 9395 -975
rect 9255 -1010 9325 -1000
rect 9255 -1040 9265 -1010
rect 9295 -1040 9325 -1010
rect 9365 -1040 9395 -1000
rect 9255 -1070 9395 -1040
rect 9255 -1100 9265 -1070
rect 9295 -1080 9395 -1070
rect 9295 -1100 9325 -1080
rect 9255 -1120 9325 -1100
rect 9365 -1120 9395 -1080
rect 9255 -1130 9395 -1120
rect 9255 -1160 9265 -1130
rect 9295 -1160 9395 -1130
rect 9255 -1175 9395 -1160
rect 1180 -1550 1380 -1540
rect 1180 -1580 1195 -1550
rect 1225 -1580 1255 -1550
rect 1285 -1580 1315 -1550
rect 1345 -1580 1380 -1550
rect 1180 -1610 1380 -1580
rect 1180 -1640 1195 -1610
rect 1225 -1640 1255 -1610
rect 1285 -1640 1315 -1610
rect 1345 -1640 1380 -1610
rect 1180 -1670 1380 -1640
rect 1180 -1710 1190 -1670
rect 1230 -1710 1270 -1670
rect 1310 -1710 1380 -1670
rect 1180 -1740 1380 -1710
rect 6580 -1785 6710 -1770
rect 6580 -1790 6650 -1785
rect 6580 -1820 6585 -1790
rect 6615 -1820 6650 -1790
rect 6580 -1825 6650 -1820
rect 6690 -1825 6710 -1785
rect 6580 -1850 6710 -1825
rect 6580 -1880 6585 -1850
rect 6615 -1880 6710 -1850
rect 6580 -1905 6710 -1880
rect 6580 -1945 6650 -1905
rect 6690 -1945 6710 -1905
rect 6580 -1970 6710 -1945
rect -1160 -2110 -960 -2095
rect -1160 -2150 -1145 -2110
rect -1105 -2150 -1020 -2110
rect -980 -2150 -960 -2110
rect -1160 -2185 -960 -2150
rect -1160 -2225 -1145 -2185
rect -1105 -2225 -1020 -2185
rect -980 -2225 -960 -2185
rect -1160 -2245 -960 -2225
rect -1160 -2275 -1140 -2245
rect -1110 -2275 -1015 -2245
rect -985 -2275 -960 -2245
rect -1160 -2295 -960 -2275
rect -740 -2750 -540 -2735
rect -740 -2780 -725 -2750
rect -695 -2780 -665 -2750
rect -635 -2780 -605 -2750
rect -575 -2780 -540 -2750
rect -740 -2815 -540 -2780
rect -740 -2855 -715 -2815
rect -675 -2855 -615 -2815
rect -575 -2855 -540 -2815
rect -740 -2885 -540 -2855
rect -740 -2925 -715 -2885
rect -675 -2925 -615 -2885
rect -575 -2925 -540 -2885
rect -740 -2935 -540 -2925
rect 9255 -3505 9380 -3470
rect -980 -3545 -740 -3530
rect -980 -3575 -965 -3545
rect -935 -3575 -905 -3545
rect -875 -3575 -845 -3545
rect -815 -3575 -785 -3545
rect -755 -3575 -740 -3545
rect -980 -3605 -740 -3575
rect -980 -3645 -965 -3605
rect -925 -3645 -885 -3605
rect -845 -3645 -805 -3605
rect -765 -3645 -740 -3605
rect -980 -3660 -740 -3645
rect 9255 -3535 9265 -3505
rect 9295 -3535 9380 -3505
rect 9255 -3565 9325 -3535
rect 9255 -3595 9265 -3565
rect 9295 -3575 9325 -3565
rect 9365 -3575 9380 -3535
rect 9295 -3595 9380 -3575
rect 9255 -3615 9380 -3595
rect 9255 -3625 9325 -3615
rect 9255 -3655 9265 -3625
rect 9295 -3655 9325 -3625
rect 9365 -3655 9380 -3615
rect 9255 -3670 9380 -3655
rect 6125 -4070 6325 -4060
rect 6125 -4100 6140 -4070
rect 6170 -4100 6200 -4070
rect 6230 -4100 6260 -4070
rect 6290 -4100 6325 -4070
rect 6125 -4115 6325 -4100
rect 6125 -4155 6135 -4115
rect 6175 -4155 6255 -4115
rect 6295 -4155 6325 -4115
rect 6125 -4160 6325 -4155
rect -820 -4585 -620 -4575
rect -820 -4615 -805 -4585
rect -775 -4615 -745 -4585
rect -715 -4615 -685 -4585
rect -655 -4615 -620 -4585
rect -820 -4630 -620 -4615
rect -820 -4670 -805 -4630
rect -765 -4670 -690 -4630
rect -650 -4670 -620 -4630
rect -820 -4685 -620 -4670
rect 290 -4580 490 -4570
rect 290 -4610 305 -4580
rect 335 -4610 365 -4580
rect 395 -4610 425 -4580
rect 455 -4610 490 -4580
rect 290 -4630 490 -4610
rect 290 -4670 305 -4630
rect 345 -4670 420 -4630
rect 460 -4670 490 -4630
rect 290 -4680 490 -4670
rect 4000 -4790 4195 -4780
rect 4000 -4820 4015 -4790
rect 4045 -4820 4075 -4790
rect 4105 -4820 4135 -4790
rect 4165 -4820 4195 -4790
rect 4000 -4845 4195 -4820
rect 4000 -4885 4020 -4845
rect 4060 -4885 4130 -4845
rect 4170 -4885 4195 -4845
rect 4000 -4900 4195 -4885
rect 8035 -4790 8230 -4780
rect 8035 -4820 8045 -4790
rect 8075 -4820 8105 -4790
rect 8135 -4820 8165 -4790
rect 8195 -4820 8230 -4790
rect 8035 -4845 8230 -4820
rect 8035 -4885 8050 -4845
rect 8090 -4885 8170 -4845
rect 8210 -4885 8230 -4845
rect 8035 -4900 8230 -4885
<< via2 >>
rect -535 4050 -495 4090
rect -415 4050 -375 4090
rect 1530 4055 1570 4095
rect 1640 4055 1680 4095
rect 5540 4055 5580 4095
rect 5655 4055 5695 4095
rect 7950 4050 7990 4090
rect 8070 4050 8110 4090
rect 7415 2355 7465 2405
rect 7415 2255 7465 2305
rect -715 440 -675 480
rect -610 440 -570 480
rect -715 370 -675 410
rect -610 370 -570 410
rect -135 435 -95 475
rect -25 435 15 475
rect -135 365 -95 405
rect -25 365 15 405
rect 465 450 505 490
rect 585 450 625 490
rect 465 370 505 410
rect 585 370 625 410
rect 9325 -1040 9365 -1000
rect 9325 -1120 9365 -1080
rect 1190 -1710 1230 -1670
rect 1270 -1710 1310 -1670
rect 6650 -1825 6690 -1785
rect 6650 -1945 6690 -1905
rect -1145 -2150 -1105 -2110
rect -1020 -2150 -980 -2110
rect -1145 -2225 -1105 -2185
rect -1020 -2225 -980 -2185
rect -715 -2855 -675 -2815
rect -615 -2855 -575 -2815
rect -715 -2925 -675 -2885
rect -615 -2925 -575 -2885
rect -965 -3645 -925 -3605
rect -885 -3645 -845 -3605
rect -805 -3645 -765 -3605
rect 9325 -3575 9365 -3535
rect 9325 -3655 9365 -3615
rect 6135 -4155 6175 -4115
rect 6255 -4155 6295 -4115
rect -805 -4670 -765 -4630
rect -690 -4670 -650 -4630
rect 305 -4670 345 -4630
rect 420 -4670 460 -4630
rect 4020 -4885 4060 -4845
rect 4130 -4885 4170 -4845
rect 8050 -4885 8090 -4845
rect 8170 -4885 8210 -4845
<< metal3 >>
rect -3162 5870 11050 5950
rect -3162 5820 -3120 5870
rect -3070 5820 -3020 5870
rect -2970 5865 7960 5870
rect -2970 5820 -535 5865
rect -3162 5815 -535 5820
rect -485 5815 -435 5865
rect -385 5815 1530 5865
rect 1580 5815 1630 5865
rect 1680 5815 5540 5865
rect 5590 5815 5640 5865
rect 5690 5820 7960 5865
rect 8010 5820 8060 5870
rect 8110 5865 11050 5870
rect 8110 5820 10810 5865
rect 5690 5815 10810 5820
rect 10860 5815 10910 5865
rect 10960 5815 11050 5865
rect -3162 5770 11050 5815
rect -3162 5720 -3120 5770
rect -3070 5720 -3020 5770
rect -2970 5765 7960 5770
rect -2970 5720 -535 5765
rect -3162 5715 -535 5720
rect -485 5715 -435 5765
rect -385 5715 1530 5765
rect 1580 5715 1630 5765
rect 1680 5715 5540 5765
rect 5590 5715 5640 5765
rect 5690 5720 7960 5765
rect 8010 5720 8060 5770
rect 8110 5765 11050 5770
rect 8110 5720 10810 5765
rect 5690 5715 10810 5720
rect 10860 5715 10910 5765
rect 10960 5715 11050 5765
rect -3162 5678 11050 5715
rect -2074 4870 10030 4930
rect -2074 4820 -2035 4870
rect -1985 4820 -1935 4870
rect -1885 4865 10030 4870
rect -1885 4820 9850 4865
rect -2074 4815 9850 4820
rect 9900 4815 9950 4865
rect 10000 4815 10030 4865
rect -2074 4770 10030 4815
rect -2074 4720 -2035 4770
rect -1985 4720 -1935 4770
rect -1885 4765 10030 4770
rect -1885 4720 9850 4765
rect -2074 4715 9850 4720
rect 9900 4715 9950 4765
rect 10000 4715 10030 4765
rect -2074 4658 10030 4715
rect 1510 4175 1710 4185
rect 1510 4125 1530 4175
rect 1580 4125 1630 4175
rect 1680 4125 1710 4175
rect -555 4100 -355 4105
rect -555 4040 -545 4100
rect -485 4040 -425 4100
rect -365 4040 -355 4100
rect -555 4035 -355 4040
rect 1510 4095 1710 4125
rect 1510 4055 1530 4095
rect 1570 4055 1640 4095
rect 1680 4055 1710 4095
rect 1510 4035 1710 4055
rect 5520 4175 5720 4185
rect 5520 4125 5540 4175
rect 5590 4125 5640 4175
rect 5690 4125 5720 4175
rect 5520 4095 5720 4125
rect 5520 4055 5540 4095
rect 5580 4055 5655 4095
rect 5695 4055 5720 4095
rect 5520 4035 5720 4055
rect 7935 4165 8135 4175
rect 7935 4115 7950 4165
rect 8000 4115 8065 4165
rect 8115 4115 8135 4165
rect 7935 4090 8135 4115
rect 7935 4050 7950 4090
rect 7990 4050 8070 4090
rect 8110 4050 8135 4090
rect 7935 4035 8135 4050
rect 7340 2405 10025 2435
rect 7340 2355 7415 2405
rect 7465 2355 9850 2405
rect 9900 2355 9950 2405
rect 10000 2355 10025 2405
rect 7340 2305 10025 2355
rect 7340 2255 7415 2305
rect 7465 2255 9850 2305
rect 9900 2255 9950 2305
rect 10000 2255 10025 2305
rect 7340 2235 10025 2255
rect -3145 525 645 555
rect -3145 475 -3125 525
rect -3075 475 -3025 525
rect -2975 490 645 525
rect -2975 480 465 490
rect -2975 475 -715 480
rect -3145 440 -715 475
rect -675 440 -610 480
rect -570 475 465 480
rect -570 440 -135 475
rect -3145 435 -135 440
rect -95 435 -25 475
rect 15 450 465 475
rect 505 450 585 490
rect 625 450 645 490
rect 15 435 645 450
rect -3145 425 645 435
rect -3145 375 -3125 425
rect -3075 375 -3025 425
rect -2975 410 645 425
rect -2975 375 -715 410
rect -3145 370 -715 375
rect -675 370 -610 410
rect -570 405 465 410
rect -570 370 -135 405
rect -3145 365 -135 370
rect -95 365 -25 405
rect 15 370 465 405
rect 505 370 585 410
rect 625 370 645 410
rect 15 365 645 370
rect -3145 355 645 365
rect 9255 -1000 10025 -975
rect 9255 -1040 9325 -1000
rect 9365 -1040 9855 -1000
rect 9255 -1050 9855 -1040
rect 9905 -1050 9955 -1000
rect 10005 -1050 10025 -1000
rect 9255 -1080 10025 -1050
rect 9255 -1120 9325 -1080
rect 9365 -1100 10025 -1080
rect 9365 -1120 9855 -1100
rect 9255 -1150 9855 -1120
rect 9905 -1150 9955 -1100
rect 10005 -1150 10025 -1100
rect 9255 -1175 10025 -1150
rect -2065 -1560 1380 -1540
rect -2065 -1610 -2035 -1560
rect -1985 -1610 -1935 -1560
rect -1885 -1610 1380 -1560
rect -2065 -1660 1380 -1610
rect -2065 -1710 -2035 -1660
rect -1985 -1710 -1935 -1660
rect -1885 -1670 1380 -1660
rect -1885 -1710 1190 -1670
rect 1230 -1710 1270 -1670
rect 1310 -1710 1380 -1670
rect -2065 -1740 1380 -1710
rect 6580 -1785 10990 -1770
rect 6580 -1825 6650 -1785
rect 6690 -1790 10990 -1785
rect 6690 -1825 10815 -1790
rect 6580 -1840 10815 -1825
rect 10865 -1840 10915 -1790
rect 10965 -1840 10990 -1790
rect 6580 -1890 10990 -1840
rect 6580 -1905 10815 -1890
rect 6580 -1945 6650 -1905
rect 6690 -1940 10815 -1905
rect 10865 -1940 10915 -1890
rect 10965 -1940 10990 -1890
rect 6690 -1945 10990 -1940
rect 6580 -1970 10990 -1945
rect -3145 -2110 -960 -2095
rect -3145 -2115 -1145 -2110
rect -3145 -2165 -3120 -2115
rect -3070 -2165 -3020 -2115
rect -2970 -2150 -1145 -2115
rect -1105 -2150 -1020 -2110
rect -980 -2150 -960 -2110
rect -2970 -2165 -960 -2150
rect -3145 -2185 -960 -2165
rect -3145 -2215 -1145 -2185
rect -3145 -2265 -3120 -2215
rect -3070 -2265 -3020 -2215
rect -2970 -2225 -1145 -2215
rect -1105 -2225 -1020 -2185
rect -980 -2225 -960 -2185
rect -2970 -2265 -960 -2225
rect -3145 -2295 -960 -2265
rect -2065 -2760 1015 -2735
rect -2065 -2810 -2045 -2760
rect -1995 -2810 -1945 -2760
rect -1895 -2810 1015 -2760
rect -2065 -2815 1015 -2810
rect -2065 -2855 -715 -2815
rect -675 -2855 -615 -2815
rect -575 -2855 1015 -2815
rect -2065 -2860 1015 -2855
rect -2065 -2910 -2045 -2860
rect -1995 -2910 -1945 -2860
rect -1895 -2885 1015 -2860
rect -1895 -2910 -715 -2885
rect -2065 -2925 -715 -2910
rect -675 -2925 -615 -2885
rect -575 -2925 1015 -2885
rect -2065 -2935 1015 -2925
rect 9255 -3495 10025 -3470
rect -2065 -3540 -740 -3515
rect -2065 -3590 -2045 -3540
rect -1995 -3590 -1945 -3540
rect -1895 -3590 -740 -3540
rect -2065 -3605 -740 -3590
rect -2065 -3640 -965 -3605
rect -2065 -3690 -2045 -3640
rect -1995 -3690 -1945 -3640
rect -1895 -3645 -965 -3640
rect -925 -3645 -885 -3605
rect -845 -3645 -805 -3605
rect -765 -3645 -740 -3605
rect -1895 -3660 -740 -3645
rect 9255 -3535 9850 -3495
rect 9255 -3575 9325 -3535
rect 9365 -3545 9850 -3535
rect 9900 -3545 9950 -3495
rect 10000 -3545 10025 -3495
rect 9365 -3575 10025 -3545
rect 9255 -3595 10025 -3575
rect 9255 -3615 9850 -3595
rect 9255 -3655 9325 -3615
rect 9365 -3645 9850 -3615
rect 9900 -3645 9950 -3595
rect 10000 -3645 10025 -3595
rect 9365 -3655 10025 -3645
rect -1895 -3690 -1865 -3660
rect 9255 -3670 10025 -3655
rect -2065 -3715 -1865 -3690
rect 6125 -4115 6325 -4110
rect 6125 -4155 6135 -4115
rect 6175 -4155 6255 -4115
rect 6295 -4155 6325 -4115
rect 6125 -4165 6325 -4155
rect 6125 -4215 6140 -4165
rect 6190 -4215 6240 -4165
rect 6290 -4215 6325 -4165
rect 6125 -4220 6325 -4215
rect -820 -4630 -620 -4620
rect -820 -4670 -805 -4630
rect -765 -4670 -690 -4630
rect -650 -4670 -620 -4630
rect -820 -4690 -620 -4670
rect -820 -4740 -805 -4690
rect -755 -4740 -705 -4690
rect -655 -4740 -620 -4690
rect 290 -4630 490 -4620
rect 290 -4670 305 -4630
rect 345 -4670 420 -4630
rect 460 -4670 490 -4630
rect 290 -4685 490 -4670
rect 290 -4735 300 -4685
rect 350 -4735 400 -4685
rect 450 -4735 490 -4685
rect 290 -4740 490 -4735
rect -820 -4750 -620 -4740
rect 4000 -4845 4195 -4830
rect 4000 -4885 4020 -4845
rect 4060 -4885 4130 -4845
rect 4170 -4885 4195 -4845
rect 4000 -4900 4195 -4885
rect 4000 -4950 4015 -4900
rect 4065 -4950 4125 -4900
rect 4175 -4950 4195 -4900
rect 4000 -4955 4195 -4950
rect 8035 -4845 8230 -4830
rect 8035 -4885 8050 -4845
rect 8090 -4885 8170 -4845
rect 8210 -4885 8230 -4845
rect 8035 -4910 8230 -4885
rect 8035 -4960 8055 -4910
rect 8105 -4960 8155 -4910
rect 8205 -4960 8230 -4910
rect 8035 -4970 8230 -4960
rect -2074 -5755 10030 -5678
rect -2074 -5805 -2035 -5755
rect -1985 -5805 -1935 -5755
rect -1885 -5760 10030 -5755
rect -1885 -5805 4020 -5760
rect -2074 -5810 4020 -5805
rect 4070 -5810 4120 -5760
rect 4170 -5810 8060 -5760
rect 8110 -5810 8160 -5760
rect 8210 -5765 10030 -5760
rect 8210 -5810 9845 -5765
rect -2074 -5815 9845 -5810
rect 9895 -5815 9945 -5765
rect 9995 -5815 10030 -5765
rect -2074 -5855 10030 -5815
rect -2074 -5905 -2035 -5855
rect -1985 -5905 -1935 -5855
rect -1885 -5860 10030 -5855
rect -1885 -5905 4020 -5860
rect -2074 -5910 4020 -5905
rect 4070 -5910 4120 -5860
rect 4170 -5910 8060 -5860
rect 8110 -5910 8160 -5860
rect 8210 -5865 10030 -5860
rect 8210 -5910 9845 -5865
rect -2074 -5915 9845 -5910
rect 9895 -5915 9945 -5865
rect 9995 -5915 10030 -5865
rect -2074 -5950 10030 -5915
rect -3162 -6855 11050 -6766
rect -3162 -6860 315 -6855
rect -3162 -6910 -3120 -6860
rect -3070 -6910 -3020 -6860
rect -2970 -6865 315 -6860
rect -2970 -6910 -800 -6865
rect -3162 -6915 -800 -6910
rect -750 -6915 -700 -6865
rect -650 -6905 315 -6865
rect 365 -6905 415 -6855
rect 465 -6905 6150 -6855
rect 6200 -6905 6250 -6855
rect 6300 -6865 11050 -6855
rect 6300 -6905 10810 -6865
rect -650 -6915 10810 -6905
rect 10860 -6915 10910 -6865
rect 10960 -6915 11050 -6865
rect -3162 -6955 11050 -6915
rect -3162 -6960 315 -6955
rect -3162 -7010 -3120 -6960
rect -3070 -7010 -3020 -6960
rect -2970 -6965 315 -6960
rect -2970 -7010 -800 -6965
rect -3162 -7015 -800 -7010
rect -750 -7015 -700 -6965
rect -650 -7005 315 -6965
rect 365 -7005 415 -6955
rect 465 -7005 6150 -6955
rect 6200 -7005 6250 -6955
rect 6300 -6965 11050 -6955
rect 6300 -7005 10810 -6965
rect -650 -7015 10810 -7005
rect 10860 -7015 10910 -6965
rect 10960 -7015 11050 -6965
rect -3162 -7038 11050 -7015
<< via3 >>
rect -3120 5820 -3070 5870
rect -3020 5820 -2970 5870
rect -535 5815 -485 5865
rect -435 5815 -385 5865
rect 1530 5815 1580 5865
rect 1630 5815 1680 5865
rect 5540 5815 5590 5865
rect 5640 5815 5690 5865
rect 7960 5820 8010 5870
rect 8060 5820 8110 5870
rect 10810 5815 10860 5865
rect 10910 5815 10960 5865
rect -3120 5720 -3070 5770
rect -3020 5720 -2970 5770
rect -535 5715 -485 5765
rect -435 5715 -385 5765
rect 1530 5715 1580 5765
rect 1630 5715 1680 5765
rect 5540 5715 5590 5765
rect 5640 5715 5690 5765
rect 7960 5720 8010 5770
rect 8060 5720 8110 5770
rect 10810 5715 10860 5765
rect 10910 5715 10960 5765
rect -2035 4820 -1985 4870
rect -1935 4820 -1885 4870
rect 9850 4815 9900 4865
rect 9950 4815 10000 4865
rect -2035 4720 -1985 4770
rect -1935 4720 -1885 4770
rect 9850 4715 9900 4765
rect 9950 4715 10000 4765
rect 1530 4125 1580 4175
rect 1630 4125 1680 4175
rect -545 4090 -485 4100
rect -545 4050 -535 4090
rect -535 4050 -495 4090
rect -495 4050 -485 4090
rect -545 4040 -485 4050
rect -425 4090 -365 4100
rect -425 4050 -415 4090
rect -415 4050 -375 4090
rect -375 4050 -365 4090
rect -425 4040 -365 4050
rect 5540 4125 5590 4175
rect 5640 4125 5690 4175
rect 7950 4115 8000 4165
rect 8065 4115 8115 4165
rect 9850 2355 9900 2405
rect 9950 2355 10000 2405
rect 9850 2255 9900 2305
rect 9950 2255 10000 2305
rect -3125 475 -3075 525
rect -3025 475 -2975 525
rect -3125 375 -3075 425
rect -3025 375 -2975 425
rect 9855 -1050 9905 -1000
rect 9955 -1050 10005 -1000
rect 9855 -1150 9905 -1100
rect 9955 -1150 10005 -1100
rect -2035 -1610 -1985 -1560
rect -1935 -1610 -1885 -1560
rect -2035 -1710 -1985 -1660
rect -1935 -1710 -1885 -1660
rect 10815 -1840 10865 -1790
rect 10915 -1840 10965 -1790
rect 10815 -1940 10865 -1890
rect 10915 -1940 10965 -1890
rect -3120 -2165 -3070 -2115
rect -3020 -2165 -2970 -2115
rect -3120 -2265 -3070 -2215
rect -3020 -2265 -2970 -2215
rect -2045 -2810 -1995 -2760
rect -1945 -2810 -1895 -2760
rect -2045 -2910 -1995 -2860
rect -1945 -2910 -1895 -2860
rect -2045 -3590 -1995 -3540
rect -1945 -3590 -1895 -3540
rect -2045 -3690 -1995 -3640
rect -1945 -3690 -1895 -3640
rect 9850 -3545 9900 -3495
rect 9950 -3545 10000 -3495
rect 9850 -3645 9900 -3595
rect 9950 -3645 10000 -3595
rect 6140 -4215 6190 -4165
rect 6240 -4215 6290 -4165
rect -805 -4740 -755 -4690
rect -705 -4740 -655 -4690
rect 300 -4735 350 -4685
rect 400 -4735 450 -4685
rect 4015 -4950 4065 -4900
rect 4125 -4950 4175 -4900
rect 8055 -4960 8105 -4910
rect 8155 -4960 8205 -4910
rect -2035 -5805 -1985 -5755
rect -1935 -5805 -1885 -5755
rect 4020 -5810 4070 -5760
rect 4120 -5810 4170 -5760
rect 8060 -5810 8110 -5760
rect 8160 -5810 8210 -5760
rect 9845 -5815 9895 -5765
rect 9945 -5815 9995 -5765
rect -2035 -5905 -1985 -5855
rect -1935 -5905 -1885 -5855
rect 4020 -5910 4070 -5860
rect 4120 -5910 4170 -5860
rect 8060 -5910 8110 -5860
rect 8160 -5910 8210 -5860
rect 9845 -5915 9895 -5865
rect 9945 -5915 9995 -5865
rect -3120 -6910 -3070 -6860
rect -3020 -6910 -2970 -6860
rect -800 -6915 -750 -6865
rect -700 -6915 -650 -6865
rect 315 -6905 365 -6855
rect 415 -6905 465 -6855
rect 6150 -6905 6200 -6855
rect 6250 -6905 6300 -6855
rect 10810 -6915 10860 -6865
rect 10910 -6915 10960 -6865
rect -3120 -7010 -3070 -6960
rect -3020 -7010 -2970 -6960
rect -800 -7015 -750 -6965
rect -700 -7015 -650 -6965
rect 315 -7005 365 -6955
rect 415 -7005 465 -6955
rect 6150 -7005 6200 -6955
rect 6250 -7005 6300 -6955
rect 10810 -7015 10860 -6965
rect 10910 -7015 10960 -6965
<< metal4 >>
rect -3162 5870 -2890 5950
rect -3162 5820 -3120 5870
rect -3070 5820 -3020 5870
rect -2970 5820 -2890 5870
rect -3162 5770 -2890 5820
rect -3162 5720 -3120 5770
rect -3070 5720 -3020 5770
rect -2970 5720 -2890 5770
rect -3162 525 -2890 5720
rect -555 5865 -355 5895
rect -555 5815 -535 5865
rect -485 5815 -435 5865
rect -385 5815 -355 5865
rect -555 5765 -355 5815
rect -555 5715 -535 5765
rect -485 5715 -435 5765
rect -385 5715 -355 5765
rect -3162 475 -3125 525
rect -3075 475 -3025 525
rect -2975 475 -2890 525
rect -3162 425 -2890 475
rect -3162 375 -3125 425
rect -3075 375 -3025 425
rect -2975 375 -2890 425
rect -3162 -2115 -2890 375
rect -3162 -2165 -3120 -2115
rect -3070 -2165 -3020 -2115
rect -2970 -2165 -2890 -2115
rect -3162 -2215 -2890 -2165
rect -3162 -2265 -3120 -2215
rect -3070 -2265 -3020 -2215
rect -2970 -2265 -2890 -2215
rect -3162 -6860 -2890 -2265
rect -2074 4870 -1802 4930
rect -2074 4820 -2035 4870
rect -1985 4820 -1935 4870
rect -1885 4820 -1802 4870
rect -2074 4770 -1802 4820
rect -2074 4720 -2035 4770
rect -1985 4720 -1935 4770
rect -1885 4720 -1802 4770
rect -2074 -1560 -1802 4720
rect -555 4100 -355 5715
rect -555 4040 -545 4100
rect -485 4040 -425 4100
rect -365 4040 -355 4100
rect -555 3995 -355 4040
rect 1510 5865 1710 5895
rect 1510 5815 1530 5865
rect 1580 5815 1630 5865
rect 1680 5815 1710 5865
rect 1510 5765 1710 5815
rect 1510 5715 1530 5765
rect 1580 5715 1630 5765
rect 1680 5715 1710 5765
rect 1510 4175 1710 5715
rect 1510 4125 1530 4175
rect 1580 4125 1630 4175
rect 1680 4125 1710 4175
rect 1510 3995 1710 4125
rect 5520 5865 5720 5895
rect 5520 5815 5540 5865
rect 5590 5815 5640 5865
rect 5690 5815 5720 5865
rect 5520 5765 5720 5815
rect 5520 5715 5540 5765
rect 5590 5715 5640 5765
rect 5690 5715 5720 5765
rect 5520 4175 5720 5715
rect 5520 4125 5540 4175
rect 5590 4125 5640 4175
rect 5690 4125 5720 4175
rect 5520 3995 5720 4125
rect 7935 5870 8135 5895
rect 7935 5820 7960 5870
rect 8010 5820 8060 5870
rect 8110 5820 8135 5870
rect 7935 5770 8135 5820
rect 7935 5720 7960 5770
rect 8010 5720 8060 5770
rect 8110 5720 8135 5770
rect 7935 4165 8135 5720
rect 10778 5865 11050 5950
rect 10778 5815 10810 5865
rect 10860 5815 10910 5865
rect 10960 5815 11050 5865
rect 10778 5765 11050 5815
rect 10778 5715 10810 5765
rect 10860 5715 10910 5765
rect 10960 5715 11050 5765
rect 7935 4115 7950 4165
rect 8000 4115 8065 4165
rect 8115 4115 8135 4165
rect 7935 3995 8135 4115
rect 9758 4865 10030 4930
rect 9758 4815 9850 4865
rect 9900 4815 9950 4865
rect 10000 4815 10030 4865
rect 9758 4765 10030 4815
rect 9758 4715 9850 4765
rect 9900 4715 9950 4765
rect 10000 4715 10030 4765
rect -2074 -1610 -2035 -1560
rect -1985 -1610 -1935 -1560
rect -1885 -1610 -1802 -1560
rect -2074 -1660 -1802 -1610
rect -2074 -1710 -2035 -1660
rect -1985 -1710 -1935 -1660
rect -1885 -1710 -1802 -1660
rect -2074 -2760 -1802 -1710
rect -2074 -2810 -2045 -2760
rect -1995 -2810 -1945 -2760
rect -1895 -2810 -1802 -2760
rect -2074 -2860 -1802 -2810
rect -2074 -2910 -2045 -2860
rect -1995 -2910 -1945 -2860
rect -1895 -2910 -1802 -2860
rect -2074 -3540 -1802 -2910
rect -2074 -3590 -2045 -3540
rect -1995 -3590 -1945 -3540
rect -1895 -3590 -1802 -3540
rect -2074 -3640 -1802 -3590
rect -2074 -3690 -2045 -3640
rect -1995 -3690 -1945 -3640
rect -1895 -3690 -1802 -3640
rect -2074 -5755 -1802 -3690
rect 9758 2405 10030 4715
rect 9758 2355 9850 2405
rect 9900 2355 9950 2405
rect 10000 2355 10030 2405
rect 9758 2305 10030 2355
rect 9758 2255 9850 2305
rect 9900 2255 9950 2305
rect 10000 2255 10030 2305
rect 9758 -1000 10030 2255
rect 9758 -1050 9855 -1000
rect 9905 -1050 9955 -1000
rect 10005 -1050 10030 -1000
rect 9758 -1100 10030 -1050
rect 9758 -1150 9855 -1100
rect 9905 -1150 9955 -1100
rect 10005 -1150 10030 -1100
rect 9758 -3495 10030 -1150
rect 9758 -3545 9850 -3495
rect 9900 -3545 9950 -3495
rect 10000 -3545 10030 -3495
rect 9758 -3595 10030 -3545
rect 9758 -3645 9850 -3595
rect 9900 -3645 9950 -3595
rect 10000 -3645 10030 -3595
rect 6125 -4165 6325 -4060
rect 6125 -4215 6140 -4165
rect 6190 -4215 6240 -4165
rect 6290 -4215 6325 -4165
rect -2074 -5805 -2035 -5755
rect -1985 -5805 -1935 -5755
rect -1885 -5805 -1802 -5755
rect -2074 -5855 -1802 -5805
rect -2074 -5905 -2035 -5855
rect -1985 -5905 -1935 -5855
rect -1885 -5905 -1802 -5855
rect -2074 -5950 -1802 -5905
rect -820 -4690 -620 -4575
rect -820 -4740 -805 -4690
rect -755 -4740 -705 -4690
rect -655 -4740 -620 -4690
rect -3162 -6910 -3120 -6860
rect -3070 -6910 -3020 -6860
rect -2970 -6910 -2890 -6860
rect -3162 -6960 -2890 -6910
rect -3162 -7010 -3120 -6960
rect -3070 -7010 -3020 -6960
rect -2970 -7010 -2890 -6960
rect -3162 -7038 -2890 -7010
rect -820 -6865 -620 -4740
rect -820 -6915 -800 -6865
rect -750 -6915 -700 -6865
rect -650 -6915 -620 -6865
rect -820 -6965 -620 -6915
rect -820 -7015 -800 -6965
rect -750 -7015 -700 -6965
rect -650 -7015 -620 -6965
rect -820 -7035 -620 -7015
rect 290 -4685 490 -4570
rect 290 -4735 300 -4685
rect 350 -4735 400 -4685
rect 450 -4735 490 -4685
rect 290 -6855 490 -4735
rect 4000 -4900 4195 -4775
rect 4000 -4950 4015 -4900
rect 4065 -4950 4125 -4900
rect 4175 -4950 4195 -4900
rect 4000 -5760 4195 -4950
rect 4000 -5810 4020 -5760
rect 4070 -5810 4120 -5760
rect 4170 -5810 4195 -5760
rect 4000 -5860 4195 -5810
rect 4000 -5910 4020 -5860
rect 4070 -5910 4120 -5860
rect 4170 -5910 4195 -5860
rect 4000 -5935 4195 -5910
rect 290 -6905 315 -6855
rect 365 -6905 415 -6855
rect 465 -6905 490 -6855
rect 290 -6955 490 -6905
rect 290 -7005 315 -6955
rect 365 -7005 415 -6955
rect 465 -7005 490 -6955
rect 290 -7035 490 -7005
rect 6125 -6855 6325 -4215
rect 8035 -4910 8230 -4780
rect 8035 -4960 8055 -4910
rect 8105 -4960 8155 -4910
rect 8205 -4960 8230 -4910
rect 8035 -5760 8230 -4960
rect 8035 -5810 8060 -5760
rect 8110 -5810 8160 -5760
rect 8210 -5810 8230 -5760
rect 8035 -5860 8230 -5810
rect 8035 -5910 8060 -5860
rect 8110 -5910 8160 -5860
rect 8210 -5910 8230 -5860
rect 8035 -5935 8230 -5910
rect 9758 -5765 10030 -3645
rect 9758 -5815 9845 -5765
rect 9895 -5815 9945 -5765
rect 9995 -5815 10030 -5765
rect 9758 -5865 10030 -5815
rect 9758 -5915 9845 -5865
rect 9895 -5915 9945 -5865
rect 9995 -5915 10030 -5865
rect 9758 -5950 10030 -5915
rect 10778 -1790 11050 5715
rect 10778 -1840 10815 -1790
rect 10865 -1840 10915 -1790
rect 10965 -1840 11050 -1790
rect 10778 -1890 11050 -1840
rect 10778 -1940 10815 -1890
rect 10865 -1940 10915 -1890
rect 10965 -1940 11050 -1890
rect 6125 -6905 6150 -6855
rect 6200 -6905 6250 -6855
rect 6300 -6905 6325 -6855
rect 6125 -6955 6325 -6905
rect 6125 -7005 6150 -6955
rect 6200 -7005 6250 -6955
rect 6300 -7005 6325 -6955
rect 6125 -7035 6325 -7005
rect 10778 -6865 11050 -1940
rect 10778 -6915 10810 -6865
rect 10860 -6915 10910 -6865
rect 10960 -6915 11050 -6865
rect 10778 -6965 11050 -6915
rect 10778 -7015 10810 -6965
rect 10860 -7015 10910 -6965
rect 10960 -7015 11050 -6965
rect 10778 -7038 11050 -7015
use ALib_DCO  ALib_DCO_0 ./../dco
timestamp 1730531556
transform 1 0 2600 0 1 -2595
box 500 -2235 6705 2990
use ALib_VCO  ALib_VCO_0 ./../vco
timestamp 1730448951
transform 1 0 -1010 0 1 520
box 0 140 10320 3515
use DLib_Quantizer  DLib_Quantizer_0 ./../quantizer
timestamp 1730532965
transform 1 0 -1105 0 1 -2315
box 95 -355 2945 365
use DLib_UpDownCounter  DLib_UpDownCounter_0 ./../count
timestamp 1730536752
transform 1 0 -570 0 1 -2993
box -440 -1577 1570 -220
use DLib_UpDownCounter  DLib_UpDownCounter_1
timestamp 1730536752
transform 1 0 -570 0 1 172
box -440 -1577 1570 -220
<< labels >>
flabel metal3 -2970 5678 -535 5950 1 FreeSans 1088 0 0 0 VDDA
port 7 nsew power input
flabel metal3 8194 4658 9758 4930 1 FreeSans 1088 0 0 0 GND
port 8 nsew ground input
<< end >>
