* NGSPICE file created from vco.ext - technology: sky130A

.subckt vco_aux_inv A VPWR VGND Y VCCA GND
X0 Y A VPWR VCCA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt vco_main_inv A VDDA VGND Y GND
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt cc_inv inp inn outp outn VDDA GND VGND
Xvco_aux_inv_0 outp VDDA VGND outn VDDA GND vco_aux_inv
Xvco_aux_inv_1 outn VDDA VGND outp VDDA GND vco_aux_inv
Xvco_main_inv_0 inp VDDA VGND outp GND vco_main_inv
Xvco_main_inv_1 inn VDDA VGND outn GND vco_main_inv
.ends

.subckt vco_ring_osc pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VGND VDDA
+ GND
Xcc_inv_0 p[4] pn[4] p[0] pn[0] VDDA GND VGND cc_inv
Xcc_inv_1 p[0] pn[0] p[1] pn[1] VDDA GND VGND cc_inv
Xcc_inv_2 p[1] pn[1] p[2] pn[2] VDDA GND VGND cc_inv
Xcc_inv_3 p[3] pn[3] p[4] pn[4] VDDA GND VGND cc_inv
Xcc_inv_4 p[2] pn[2] p[3] pn[3] VDDA GND VGND cc_inv
.ends

.subckt sky130_fd_pr__res_generic_po_DKCPUZ a_n48_200# a_n48_n630#
R0 a_n48_200# a_n48_n630# sky130_fd_pr__res_generic_po w=0.48 l=2
.ends


.subckt vco VCCD ENB p[4] Anlg_in VCCA VPWR GND
Xvco_ring_osc_0 vco_ring_osc_0/pn[0] vco_ring_osc_0/pn[1] vco_ring_osc_0/pn[2] vco_ring_osc_0/pn[3]
+ vco_ring_osc_0/pn[4] vco_ring_osc_0/p[0] vco_ring_osc_0/p[1] vco_ring_osc_0/p[2]
+ vco_ring_osc_0/p[3] p[4] vco_ring_osc_0/VGND VPWR GND vco_ring_osc
Xsky130_fd_pr__res_generic_po_DKCPUZ_0 Anlg_in vco_ring_osc_0/VGND sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_pr__res_generic_po_DKCPUZ_1 vco_ring_osc_0/VGND GND sky130_fd_pr__res_generic_po_DKCPUZ
Xsky130_fd_sc_hd__einvp_1_0 VCCD ENB GND GND VCCD VCCD vco_ring_osc_0/pn[4] sky130_fd_sc_hd__einvp_1
.ends


