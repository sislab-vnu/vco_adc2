magic
tech sky130A
timestamp 1725081791
<< nwell >>
rect 1425 500 1465 540
rect 1830 -40 1890 540
<< poly >>
rect 1060 -45 1425 -40
rect 1060 -65 1150 -45
rect 1170 -65 1190 -45
rect 1210 -65 1230 -45
rect 1250 -65 1425 -45
rect 1465 -45 1830 -40
rect 1465 -65 1520 -45
rect 1540 -65 1560 -45
rect 1580 -65 1600 -45
rect 1620 -65 1830 -45
<< polycont >>
rect 1150 -65 1170 -45
rect 1190 -65 1210 -45
rect 1230 -65 1250 -45
rect 1520 -65 1540 -45
rect 1560 -65 1580 -45
rect 1600 -65 1620 -45
<< locali >>
rect 1020 590 1870 630
rect 1020 500 1060 590
rect 1830 500 1870 590
rect 1140 -45 1260 -20
rect 1140 -65 1150 -45
rect 1170 -65 1190 -45
rect 1210 -65 1230 -45
rect 1250 -65 1260 -45
rect 1140 -85 1260 -65
rect 1425 -105 1465 0
rect 1510 -45 1630 -20
rect 1510 -65 1520 -45
rect 1540 -65 1560 -45
rect 1580 -65 1600 -45
rect 1620 -65 1630 -45
rect 1510 -85 1630 -65
rect 1020 -595 1060 -505
rect 1830 -595 1870 -505
rect 1020 -635 1870 -595
<< viali >>
rect 1150 -65 1170 -45
rect 1190 -65 1210 -45
rect 1230 -65 1250 -45
rect 1520 -65 1540 -45
rect 1560 -65 1580 -45
rect 1600 -65 1620 -45
<< metal1 >>
rect 1140 -45 1630 -20
rect 1140 -65 1150 -45
rect 1170 -65 1190 -45
rect 1210 -65 1230 -45
rect 1250 -65 1520 -45
rect 1540 -65 1560 -45
rect 1580 -65 1600 -45
rect 1620 -65 1630 -45
rect 1140 -85 1630 -65
use nmos_vco  nmos_vco_0
timestamp 1724742977
transform 1 0 1060 0 1 -505
box -60 -130 830 490
use pmos_vco  pmos_vco_0
timestamp 1725081437
transform 1 0 1060 0 1 0
box -60 -90 830 630
<< labels >>
rlabel locali 1445 -5 1445 -5 1 D
port 1 n
rlabel metal1 1445 -50 1445 -50 1 G
port 2 n
rlabel locali 1440 600 1440 600 1 S_P
port 3 n
rlabel locali 1445 -600 1445 -600 1 S_N
port 4 n
rlabel nwell 1445 530 1445 530 1 VPWR
port 5 n
<< end >>
