magic
tech sky130A
timestamp 1730448951
<< nwell >>
rect 2765 1450 2885 1610
<< pwell >>
rect 2775 1330 2885 1420
<< psubdiff >>
rect 2820 1390 2860 1405
rect 2820 1370 2830 1390
rect 2850 1370 2860 1390
rect 2820 1355 2860 1370
<< nsubdiff >>
rect 2820 1540 2860 1555
rect 2820 1520 2830 1540
rect 2850 1520 2860 1540
rect 2820 1505 2860 1520
<< psubdiffcont >>
rect 2830 1370 2850 1390
<< nsubdiffcont >>
rect 2830 1520 2850 1540
<< locali >>
rect 390 3475 830 3515
rect 2695 1945 2735 1950
rect 2695 1905 3425 1945
rect 2695 1900 2735 1905
rect 3425 1740 3520 1800
rect 2820 1540 2860 1555
rect 2820 1520 2830 1540
rect 2850 1520 2860 1540
rect 2820 1505 2860 1520
rect 2495 1455 2575 1485
rect 2780 1475 2805 1485
rect 2790 1455 2805 1475
rect 2780 1435 2805 1455
rect 2925 1475 2975 1485
rect 2925 1445 2935 1475
rect 2965 1445 2975 1475
rect 2820 1390 2860 1405
rect 2820 1370 2830 1390
rect 2850 1370 2860 1390
rect 2820 1355 2860 1370
rect 2925 190 2975 1445
rect 2925 140 3360 190
<< viali >>
rect 2830 1520 2850 1540
rect 2770 1455 2790 1475
rect 2935 1445 2965 1475
rect 2755 1370 2772 1387
rect 2830 1370 2850 1390
<< metal1 >>
rect 2045 1895 2085 1950
rect 2555 1685 2975 1735
rect 2565 1615 2615 1685
rect 2820 1540 2860 1685
rect 2820 1520 2830 1540
rect 2850 1520 2860 1540
rect 2820 1505 2860 1520
rect 2745 1475 2805 1495
rect 2745 1455 2770 1475
rect 2790 1465 2805 1475
rect 2925 1475 2975 1685
rect 2925 1465 2935 1475
rect 2790 1455 2935 1465
rect 2745 1445 2935 1455
rect 2965 1445 2975 1475
rect 2745 1435 2975 1445
rect 2740 1400 2785 1410
rect 2445 1387 2785 1400
rect 2445 1370 2755 1387
rect 2772 1370 2785 1387
rect 2445 1115 2495 1370
rect 2740 1365 2785 1370
rect 2820 1390 2860 1405
rect 3115 1390 3165 2100
rect 4200 1795 4250 1860
rect 4115 1740 4250 1795
rect 4200 1710 4250 1740
rect 2820 1370 2830 1390
rect 2850 1370 3165 1390
rect 2820 1360 3165 1370
rect 2820 1355 2860 1360
rect 3115 1325 3165 1360
rect 2785 1295 3165 1325
rect 2955 1075 3300 1125
rect 2970 440 3320 490
use sky130_fd_pr__res_generic_po_DKCPUZ  sky130_fd_pr__res_generic_po_DKCPUZ_0
timestamp 1725958087
transform 0 -1 2390 1 0 1924
box -24 -315 24 315
use sky130_fd_pr__res_generic_po_DKCPUZ  sky130_fd_pr__res_generic_po_DKCPUZ_1
timestamp 1725958087
transform 0 -1 3820 1 0 1769
box -24 -315 24 315
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 2564 0 1 1319
box -19 -24 249 296
use x5s_cc_osc  x5s_cc_osc_0
timestamp 1730447269
transform 1 0 300 0 1 2100
box -300 -1950 10020 1415
<< labels >>
rlabel metal1 2055 1950 2055 1950 1 Anlg_in
port 1 n
rlabel locali 2510 1485 2510 1485 1 ENB
port 2 n
rlabel metal1 3065 490 3065 490 1 p[4]
port 3 n
rlabel locali 575 3515 575 3515 1 VDDA
port 4 n
rlabel metal1 4180 1795 4180 1795 1 GND
port 5 n
rlabel metal1 3155 1125 3155 1125 1 pn[4]
rlabel locali 3360 1945 3360 1945 1 Vctrl
<< end >>
