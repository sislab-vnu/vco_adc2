magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect 750 1970 790 2010
rect -90 1850 260 1950
rect 3290 1810 3730 2050
rect 3800 1850 3810 1950
rect 4830 1650 4870 1690
rect 4830 1570 4870 1610
<< poly >>
rect 2150 1177 2190 1180
rect 2150 1143 2153 1177
rect 2187 1143 2190 1177
rect 2150 1140 2190 1143
rect 2230 1177 2270 1180
rect 2230 1143 2233 1177
rect 2267 1143 2270 1177
rect 2230 1140 2270 1143
rect 2310 1177 2350 1180
rect 2310 1143 2313 1177
rect 2347 1143 2350 1177
rect 2310 1140 2350 1143
rect 3120 1177 3160 1180
rect 3120 1143 3123 1177
rect 3157 1143 3160 1177
rect 3120 1140 3160 1143
rect 3200 1177 3240 1180
rect 3200 1143 3203 1177
rect 3237 1143 3240 1177
rect 3200 1140 3240 1143
rect 3280 1177 3320 1180
rect 3280 1143 3283 1177
rect 3317 1143 3320 1177
rect 3280 1140 3320 1143
<< polycont >>
rect 2153 1143 2187 1177
rect 2233 1143 2267 1177
rect 2313 1143 2347 1177
rect 3123 1143 3157 1177
rect 3203 1143 3237 1177
rect 3283 1143 3317 1177
<< locali >>
rect 1610 2450 4190 2530
rect 1820 2270 1900 2450
rect 2910 2270 2990 2450
rect 750 2007 790 2010
rect 750 1973 753 2007
rect 787 1973 790 2007
rect 750 1970 790 1973
rect 3740 2007 3780 2010
rect 3740 1973 3743 2007
rect 3777 1973 3780 2007
rect 3740 1970 3780 1973
rect 750 1927 790 1930
rect 750 1893 753 1927
rect 787 1893 790 1927
rect 750 1890 790 1893
rect 3740 1927 3780 1930
rect 3740 1893 3743 1927
rect 3777 1893 3780 1927
rect 3740 1890 3780 1893
rect 750 1847 790 1850
rect 750 1813 753 1847
rect 787 1813 790 1847
rect 750 1810 790 1813
rect 3740 1847 3780 1850
rect 3740 1813 3743 1847
rect 3777 1813 3780 1847
rect 3740 1810 3780 1813
rect 2650 1687 2690 1690
rect 2650 1653 2653 1687
rect 2687 1653 2690 1687
rect 2650 1650 2690 1653
rect 4830 1687 4870 1690
rect 4830 1653 4833 1687
rect 4867 1653 4870 1687
rect 4830 1650 4870 1653
rect 2650 1607 2690 1610
rect 2650 1573 2653 1607
rect 2687 1573 2690 1607
rect 2650 1570 2690 1573
rect 4830 1607 4870 1610
rect 4830 1573 4833 1607
rect 4867 1573 4870 1607
rect 4830 1570 4870 1573
rect 2650 1527 2690 1530
rect 2650 1493 2653 1527
rect 2687 1493 2690 1527
rect 2650 1490 2690 1493
rect 4830 1527 4870 1530
rect 4830 1493 4833 1527
rect 4867 1493 4870 1527
rect 4830 1490 4870 1493
rect 2130 1210 2370 1230
rect 3100 1220 3340 1230
rect 1300 1177 2370 1210
rect 1300 1143 2153 1177
rect 2187 1143 2233 1177
rect 2267 1143 2313 1177
rect 2347 1143 2370 1177
rect 1300 1110 2370 1143
rect 2710 1177 3340 1220
rect 2710 1143 3123 1177
rect 3157 1143 3203 1177
rect 3237 1143 3283 1177
rect 3317 1143 3340 1177
rect 2710 1120 3340 1143
rect 1300 990 1400 1110
rect 2130 1100 2370 1110
rect 3100 1100 3340 1120
rect 810 890 1400 990
rect 4830 717 4870 720
rect 4830 683 4833 717
rect 4867 683 4870 717
rect 4830 680 4870 683
rect 4830 637 4870 640
rect 4830 603 4833 637
rect 4867 603 4870 637
rect 4830 600 4870 603
rect 4830 557 4870 560
rect 4830 523 4833 557
rect 4867 523 4870 557
rect 4830 520 4870 523
rect 1820 80 1900 260
rect 2910 80 2990 260
rect 1620 0 4000 80
<< viali >>
rect 753 1973 787 2007
rect 3743 1973 3777 2007
rect 753 1893 787 1927
rect 3743 1893 3777 1927
rect 753 1813 787 1847
rect 3743 1813 3777 1847
rect 2653 1653 2687 1687
rect 4833 1653 4867 1687
rect 2653 1573 2687 1607
rect 4833 1573 4867 1607
rect 2653 1493 2687 1527
rect 4833 1493 4867 1527
rect 2153 1143 2187 1177
rect 2233 1143 2267 1177
rect 2313 1143 2347 1177
rect 3123 1143 3157 1177
rect 3203 1143 3237 1177
rect 3283 1143 3317 1177
rect 4833 683 4867 717
rect 4833 603 4867 637
rect 4833 523 4867 557
<< metal1 >>
rect -220 2730 3940 2830
rect -220 2280 -140 2730
rect 1680 2280 1760 2730
rect 2770 2280 2850 2730
rect 3860 2280 3940 2730
rect 730 2007 810 2050
rect 730 1973 753 2007
rect 787 1973 810 2007
rect 730 1950 810 1973
rect 3720 2007 3800 2050
rect 3720 1973 3743 2007
rect 3777 1973 3800 2007
rect 3720 1950 3800 1973
rect -260 1850 540 1950
rect 440 1230 540 1850
rect 730 1927 5740 1950
rect 730 1893 753 1927
rect 787 1893 3743 1927
rect 3777 1893 5740 1927
rect 730 1850 5740 1893
rect 730 1847 810 1850
rect 730 1813 753 1847
rect 787 1813 810 1847
rect 730 1770 810 1813
rect 2200 1230 2300 1850
rect 3720 1847 3800 1850
rect 3720 1813 3743 1847
rect 3777 1813 3800 1847
rect 3720 1770 3800 1813
rect 2630 1687 2710 1710
rect 2630 1653 2653 1687
rect 2687 1653 2710 1687
rect 2630 1640 2710 1653
rect 4810 1687 4890 1710
rect 4810 1653 4833 1687
rect 4867 1653 4890 1687
rect 4810 1640 4890 1653
rect 2630 1607 4890 1640
rect 2630 1573 2653 1607
rect 2687 1573 4833 1607
rect 4867 1573 4890 1607
rect 2630 1540 4890 1573
rect 2630 1527 2710 1540
rect 2630 1493 2653 1527
rect 2687 1493 2710 1527
rect 2630 1470 2710 1493
rect 3170 1230 3270 1540
rect 4810 1527 4890 1540
rect 4810 1493 4833 1527
rect 4867 1493 4890 1527
rect 4810 1470 4890 1493
rect 2130 1177 2370 1230
rect 2130 1143 2153 1177
rect 2187 1143 2233 1177
rect 2267 1143 2313 1177
rect 2347 1143 2370 1177
rect 2130 1100 2370 1143
rect 3100 1177 3340 1230
rect 3100 1143 3123 1177
rect 3157 1143 3203 1177
rect 3237 1143 3283 1177
rect 3317 1143 3340 1177
rect 3100 1100 3340 1143
rect 4070 1110 4240 1210
rect 4070 680 4170 1110
rect -260 580 4170 680
rect 4810 717 4890 740
rect 4810 683 4833 717
rect 4867 683 4890 717
rect 4810 680 4890 683
rect 4810 637 5740 680
rect 4810 603 4833 637
rect 4867 603 5740 637
rect 4810 580 5740 603
rect 4810 557 4890 580
rect 4810 523 4833 557
rect 4867 523 4890 557
rect 4810 500 4890 523
rect -220 -200 -140 250
rect 1680 -200 1760 250
rect 2770 -200 2850 250
rect 3860 -200 3940 250
rect -220 -300 3940 -200
use vco_aux_inv  vco_aux_inv_0
timestamp 1729593089
transform 1 0 1900 0 1 1280
box -260 -1100 850 1070
use vco_aux_inv  vco_aux_inv_1
timestamp 1729593089
transform 1 0 2990 0 1 1280
box -260 -1100 850 1070
use vco_main_inv  vco_main_inv_0
timestamp 1729593089
transform 1 0 0 0 1 1270
box -260 -1270 1660 1260
use vco_main_inv  vco_main_inv_1
timestamp 1729593089
transform 1 0 4080 0 1 1270
box -260 -1270 1660 1260
<< labels >>
rlabel metal1 s -260 1900 -260 1900 4 inp
rlabel metal1 s -260 620 -260 620 4 inn
rlabel locali s 2830 2530 2830 2530 4 VPWR
rlabel locali s 2830 0 2830 0 4 VGND
rlabel metal1 s 5740 1900 5740 1900 4 outp
rlabel metal1 s 5740 620 5740 620 4 outn
rlabel metal1 s -180 2830 -180 2830 4 VCCA
rlabel metal1 s -190 -300 -190 -300 4 GND
<< end >>
