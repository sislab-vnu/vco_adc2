magic
tech sky130A
magscale 1 2
timestamp 1724225640
<< poly >>
rect -40 579 40 595
rect -40 545 -24 579
rect 24 545 40 579
rect -40 165 40 545
rect -40 -545 40 -165
rect -40 -579 -24 -545
rect 24 -579 40 -545
rect -40 -595 40 -579
<< polycont >>
rect -24 545 24 579
rect -24 -579 24 -545
<< npolyres >>
rect -40 -165 40 165
<< locali >>
rect -40 545 -24 579
rect 24 545 40 579
rect -40 -579 -24 -545
rect 24 -579 40 -545
<< viali >>
rect -24 545 24 579
rect -24 182 24 545
rect -24 -545 24 -182
rect -24 -579 24 -545
<< metal1 >>
rect -30 579 30 591
rect -30 182 -24 579
rect 24 182 30 579
rect -30 170 30 182
rect -30 -182 30 -170
rect -30 -579 -24 -182
rect 24 -579 30 -182
rect -30 -591 30 -579
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.397 l 1.650 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 200.327 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
