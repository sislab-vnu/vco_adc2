.title Up Down Counter
* Written for	: NGSPICE
* Lib				:	testing
* Cell name	 
* Author duck-manh-tran
******************************************************

.lib /home/dkit/efabless/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc ../library/analog_lib.spice
.inc ../library/digital_lib.spice
.global gnd vdd
.param mc_mm_switch=1
*_____________sub circuits_____________*

.subckt DL_BLK	A VGND VNB VPB VPWR Y0 Y1 Y2 Y3 Y4 Y5 	$delay 1.6 ns
X_delay0 A  VGND VNB VPB VPWR Y0 sky130_fd_sc_hd__dlygate4sd1_1
X_delay1 Y0 VGND VNB VPB VPWR Y1 sky130_fd_sc_hd__dlygate4sd2_1
X_delay2 Y1 VGND VNB VPB VPWR Y2 sky130_fd_sc_hd__dlygate4sd3_1
X_delay3 Y2 VGND VNB VPB VPWR Y3 sky130_fd_sc_hd__dlygate4sd3_1
X_delay4 Y3 VGND VNB VPB VPWR Y4 sky130_fd_sc_hd__dlygate4sd3_1
X_delay5 Y4 VGND VNB VPB VPWR Y5 sky130_fd_sc_hd__dlygate4sd3_1
.ends

.subckt ADC_DigitalLib_UDCnter UP DOWN VGND VNB VPB VPWR Dout
X0 UP   Q2_INV VGND VNB VPB VPWR Q1_D2 sky130_fd_sc_hd__dfxtp_1
X1 DOWN Q1_D2  VGND VNB VPB VPWR Q2 sky130_fd_sc_hd__dfxtp_1
X2 Q2 VGND VNB VPB VPWR Q2_INV sky130_fd_sc_hd__inv_2
X3 Q1_D2 Q2 VGND VNB VPB VPWR Dout sky130_fd_sc_hd__xor2_1
.ends


*_____________UpDown Counter testbench__________________*

* UP DOWN COUNTER
* X_UD_count up_pulse down_pulse gnd gnd vdd vdd Dout ADC_DigitalLib_UDCnter

X_inv_0  rst 	gnd gnd vdd vdd rstBi sky130_fd_sc_ms__inv_2
X_buf_0  UP 	gnd gnd vdd vdd up_buf sky130_fd_sc_ms__buf_2
X_upFF_0 UP_buf Q2N rstBi gnd gnd vdd vdd Q1 sky130_fd_sc_ms__dfrtp_1
X_buf_1  Q1 gnd gnd vdd vdd Q1_buf sky130_fd_sc_ms__buf_2
X_buf_2  DOWN gnd gnd vdd vdd dwn_buf sky130_fd_sc_ms__buf_2
X_dwLATCH_0 pseudo_Q1_buf dwn_buf xxxx gnd gnd vdd vdd Q2 sky130_fd_sc_ms__dlrtp_1
X_inv_1  Q2 gnd gnd vdd vdd Q2N sky130_fd_sc_ms__inv_2
X_xor_0  Q1_buf Q2 gnd gnd vdd vdd Dout sky130_fd_sc_ms__xor2_1
X_buf_3  Dout gnd gnd vdd vdd Dout_buf sky130_fd_sc_ms__buf_2

* Ring Oscillator
X_vco_0 ENB Anlg_in GND GND VDD VDD up Vctrl ADC_AnalogLib_VCO

* DELAY BLOCK
*X_dlblk_0 sig_pwl 0 0 VDD VDD DL1 DL2 DL3 DL4 DL5 DL6 DL_BLK

* REFERENCE VOLTAGES
V1 vdd gnd DC=1.8
V1_ vdd_osc gnd DC = 1.8
V2  Anlg_in gnd DC = 0.9
*V2 up_pulse   gnd DC=0 PULSE( 0.7 1.8 40n 10n 10n 40n 100n )
V3 down gnd DC=0 PULSE( 0 1.8 0 0.2n 0.2n 17n 41.67n )
V4 enb gnd DC=0 PULSE( 0 1.8 0 20n 20n 200n 1 ) 
V5 sig_pwl gnd DC=0 PULSE( 0 1.8 0 0.1n 0.1n 50n 200n )
V6 pseudo_Q1_buf gnd DC=0 PULSE( 0 1.8 0 0.1n 0.1n 200n 400n )

* CONTROL TESTBENCH
.control
tran 0.01n 2u
plot up_pulse down_pulse Dout 
plot Dout up_pulse down_pulse 
*plot sig_pwl DL1 DL2 DL3 DL4 DL5
.endc
