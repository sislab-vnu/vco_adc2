magic
tech sky130A
timestamp 1726019674
<< nwell >>
rect -130 -40 830 540
<< pwell >>
rect -130 -545 830 -65
<< nmos >>
rect 0 -505 365 -105
rect 405 -505 770 -105
<< pmos >>
rect 0 0 365 500
rect 405 0 770 500
<< ndiff >>
rect -40 -115 0 -105
rect -40 -135 -30 -115
rect -10 -135 0 -115
rect -40 -155 0 -135
rect -40 -175 -30 -155
rect -10 -175 0 -155
rect -40 -195 0 -175
rect -40 -215 -30 -195
rect -10 -215 0 -195
rect -40 -235 0 -215
rect -40 -255 -30 -235
rect -10 -255 0 -235
rect -40 -275 0 -255
rect -40 -295 -30 -275
rect -10 -295 0 -275
rect -40 -315 0 -295
rect -40 -335 -30 -315
rect -10 -335 0 -315
rect -40 -355 0 -335
rect -40 -375 -30 -355
rect -10 -375 0 -355
rect -40 -395 0 -375
rect -40 -415 -30 -395
rect -10 -415 0 -395
rect -40 -435 0 -415
rect -40 -455 -30 -435
rect -10 -455 0 -435
rect -40 -475 0 -455
rect -40 -495 -30 -475
rect -10 -495 0 -475
rect -40 -505 0 -495
rect 365 -115 405 -105
rect 365 -135 375 -115
rect 395 -135 405 -115
rect 365 -155 405 -135
rect 365 -175 375 -155
rect 395 -175 405 -155
rect 365 -195 405 -175
rect 365 -215 375 -195
rect 395 -215 405 -195
rect 365 -235 405 -215
rect 365 -255 375 -235
rect 395 -255 405 -235
rect 365 -275 405 -255
rect 365 -295 375 -275
rect 395 -295 405 -275
rect 365 -315 405 -295
rect 365 -335 375 -315
rect 395 -335 405 -315
rect 365 -355 405 -335
rect 365 -375 375 -355
rect 395 -375 405 -355
rect 365 -395 405 -375
rect 365 -415 375 -395
rect 395 -415 405 -395
rect 365 -435 405 -415
rect 365 -455 375 -435
rect 395 -455 405 -435
rect 365 -475 405 -455
rect 365 -495 375 -475
rect 395 -495 405 -475
rect 365 -505 405 -495
rect 770 -115 810 -105
rect 770 -135 780 -115
rect 800 -135 810 -115
rect 770 -155 810 -135
rect 770 -175 780 -155
rect 800 -175 810 -155
rect 770 -195 810 -175
rect 770 -215 780 -195
rect 800 -215 810 -195
rect 770 -235 810 -215
rect 770 -255 780 -235
rect 800 -255 810 -235
rect 770 -275 810 -255
rect 770 -295 780 -275
rect 800 -295 810 -275
rect 770 -315 810 -295
rect 770 -335 780 -315
rect 800 -335 810 -315
rect 770 -355 810 -335
rect 770 -375 780 -355
rect 800 -375 810 -355
rect 770 -395 810 -375
rect 770 -415 780 -395
rect 800 -415 810 -395
rect 770 -435 810 -415
rect 770 -455 780 -435
rect 800 -455 810 -435
rect 770 -475 810 -455
rect 770 -495 780 -475
rect 800 -495 810 -475
rect 770 -505 810 -495
<< pdiff >>
rect -40 490 0 500
rect -40 470 -30 490
rect -10 470 0 490
rect -40 450 0 470
rect -40 430 -30 450
rect -10 430 0 450
rect -40 410 0 430
rect -40 390 -30 410
rect -10 390 0 410
rect -40 370 0 390
rect -40 350 -30 370
rect -10 350 0 370
rect -40 330 0 350
rect -40 310 -30 330
rect -10 310 0 330
rect -40 290 0 310
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 365 490 405 500
rect 365 470 375 490
rect 395 470 405 490
rect 365 450 405 470
rect 365 430 375 450
rect 395 430 405 450
rect 365 410 405 430
rect 365 390 375 410
rect 395 390 405 410
rect 365 370 405 390
rect 365 350 375 370
rect 395 350 405 370
rect 365 330 405 350
rect 365 310 375 330
rect 395 310 405 330
rect 365 290 405 310
rect 365 270 375 290
rect 395 270 405 290
rect 365 250 405 270
rect 365 230 375 250
rect 395 230 405 250
rect 365 210 405 230
rect 365 190 375 210
rect 395 190 405 210
rect 365 170 405 190
rect 365 150 375 170
rect 395 150 405 170
rect 365 130 405 150
rect 365 110 375 130
rect 395 110 405 130
rect 365 90 405 110
rect 365 70 375 90
rect 395 70 405 90
rect 365 50 405 70
rect 365 30 375 50
rect 395 30 405 50
rect 365 0 405 30
rect 770 490 810 500
rect 770 470 780 490
rect 800 470 810 490
rect 770 450 810 470
rect 770 430 780 450
rect 800 430 810 450
rect 770 410 810 430
rect 770 390 780 410
rect 800 390 810 410
rect 770 370 810 390
rect 770 350 780 370
rect 800 350 810 370
rect 770 330 810 350
rect 770 310 780 330
rect 800 310 810 330
rect 770 290 810 310
rect 770 270 780 290
rect 800 270 810 290
rect 770 250 810 270
rect 770 230 780 250
rect 800 230 810 250
rect 770 210 810 230
rect 770 190 780 210
rect 800 190 810 210
rect 770 170 810 190
rect 770 150 780 170
rect 800 150 810 170
rect 770 130 810 150
rect 770 110 780 130
rect 800 110 810 130
rect 770 90 810 110
rect 770 70 780 90
rect 800 70 810 90
rect 770 50 810 70
rect 770 30 780 50
rect 800 30 810 50
rect 770 0 810 30
<< ndiffc >>
rect -30 -135 -10 -115
rect -30 -175 -10 -155
rect -30 -215 -10 -195
rect -30 -255 -10 -235
rect -30 -295 -10 -275
rect -30 -335 -10 -315
rect -30 -375 -10 -355
rect -30 -415 -10 -395
rect -30 -455 -10 -435
rect -30 -495 -10 -475
rect 375 -135 395 -115
rect 375 -175 395 -155
rect 375 -215 395 -195
rect 375 -255 395 -235
rect 375 -295 395 -275
rect 375 -335 395 -315
rect 375 -375 395 -355
rect 375 -415 395 -395
rect 375 -455 395 -435
rect 375 -495 395 -475
rect 780 -135 800 -115
rect 780 -175 800 -155
rect 780 -215 800 -195
rect 780 -255 800 -235
rect 780 -295 800 -275
rect 780 -335 800 -315
rect 780 -375 800 -355
rect 780 -415 800 -395
rect 780 -455 800 -435
rect 780 -495 800 -475
<< pdiffc >>
rect -30 470 -10 490
rect -30 430 -10 450
rect -30 390 -10 410
rect -30 350 -10 370
rect -30 310 -10 330
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 375 470 395 490
rect 375 430 395 450
rect 375 390 395 410
rect 375 350 395 370
rect 375 310 395 330
rect 375 270 395 290
rect 375 230 395 250
rect 375 190 395 210
rect 375 150 395 170
rect 375 110 395 130
rect 375 70 395 90
rect 375 30 395 50
rect 780 470 800 490
rect 780 430 800 450
rect 780 390 800 410
rect 780 350 800 370
rect 780 310 800 330
rect 780 270 800 290
rect 780 230 800 250
rect 780 190 800 210
rect 780 150 800 170
rect 780 110 800 130
rect 780 70 800 90
rect 780 30 800 50
<< psubdiff >>
rect -110 -475 -70 -460
rect -110 -495 -100 -475
rect -80 -495 -70 -475
rect -110 -510 -70 -495
<< nsubdiff >>
rect -110 490 -70 505
rect -110 470 -100 490
rect -80 470 -70 490
rect -110 455 -70 470
<< psubdiffcont >>
rect -100 -495 -80 -475
<< nsubdiffcont >>
rect -100 470 -80 490
<< poly >>
rect 0 500 365 540
rect 405 500 770 540
rect 0 -15 365 0
rect 405 -15 770 0
rect 0 -45 770 -15
rect 0 -65 90 -45
rect 110 -65 130 -45
rect 150 -65 170 -45
rect 190 -65 460 -45
rect 480 -65 500 -45
rect 520 -65 540 -45
rect 560 -65 770 -45
rect 0 -90 770 -65
rect 0 -105 365 -90
rect 405 -105 770 -90
rect 0 -545 365 -505
rect 405 -545 770 -505
<< polycont >>
rect 90 -65 110 -45
rect 130 -65 150 -45
rect 170 -65 190 -45
rect 460 -65 480 -45
rect 500 -65 520 -45
rect 540 -65 560 -45
<< locali >>
rect -40 590 810 630
rect -110 490 -70 505
rect -110 470 -100 490
rect -80 470 -70 490
rect -110 455 -70 470
rect -40 490 0 590
rect -40 470 -30 490
rect -10 470 0 490
rect -40 450 0 470
rect -40 430 -30 450
rect -10 430 0 450
rect -40 410 0 430
rect -40 390 -30 410
rect -10 390 0 410
rect -40 370 0 390
rect -40 350 -30 370
rect -10 350 0 370
rect -40 330 0 350
rect -40 310 -30 330
rect -10 310 0 330
rect -40 290 0 310
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 365 490 405 500
rect 365 470 375 490
rect 395 470 405 490
rect 365 450 405 470
rect 365 430 375 450
rect 395 430 405 450
rect 365 410 405 430
rect 365 390 375 410
rect 395 390 405 410
rect 365 370 405 390
rect 365 350 375 370
rect 395 350 405 370
rect 365 330 405 350
rect 365 310 375 330
rect 395 310 405 330
rect 365 290 405 310
rect 365 270 375 290
rect 395 270 405 290
rect 365 250 405 270
rect 365 230 375 250
rect 395 230 405 250
rect 365 210 405 230
rect 365 190 375 210
rect 395 190 405 210
rect 365 170 405 190
rect 365 150 375 170
rect 395 150 405 170
rect 365 130 405 150
rect 365 110 375 130
rect 395 110 405 130
rect 365 90 405 110
rect 365 70 375 90
rect 395 70 405 90
rect 365 50 405 70
rect 365 30 375 50
rect 395 30 405 50
rect 80 -45 200 -20
rect 80 -65 90 -45
rect 110 -65 130 -45
rect 150 -65 170 -45
rect 190 -65 200 -45
rect 80 -85 200 -65
rect -40 -115 0 -105
rect -40 -135 -30 -115
rect -10 -135 0 -115
rect -40 -155 0 -135
rect -40 -175 -30 -155
rect -10 -175 0 -155
rect -40 -195 0 -175
rect -40 -215 -30 -195
rect -10 -215 0 -195
rect -40 -235 0 -215
rect -40 -255 -30 -235
rect -10 -255 0 -235
rect -40 -275 0 -255
rect -40 -295 -30 -275
rect -10 -295 0 -275
rect -40 -315 0 -295
rect -40 -335 -30 -315
rect -10 -335 0 -315
rect -40 -355 0 -335
rect -40 -375 -30 -355
rect -10 -375 0 -355
rect -40 -395 0 -375
rect -40 -415 -30 -395
rect -10 -415 0 -395
rect -40 -435 0 -415
rect -40 -455 -30 -435
rect -10 -455 0 -435
rect -110 -475 -70 -460
rect -110 -495 -100 -475
rect -80 -495 -70 -475
rect -110 -510 -70 -495
rect -40 -475 0 -455
rect -40 -495 -30 -475
rect -10 -495 0 -475
rect -40 -595 0 -495
rect 365 -115 405 30
rect 770 490 810 590
rect 770 470 780 490
rect 800 470 810 490
rect 770 450 810 470
rect 770 430 780 450
rect 800 430 810 450
rect 770 410 810 430
rect 770 390 780 410
rect 800 390 810 410
rect 770 370 810 390
rect 770 350 780 370
rect 800 350 810 370
rect 770 330 810 350
rect 770 310 780 330
rect 800 310 810 330
rect 770 290 810 310
rect 770 270 780 290
rect 800 270 810 290
rect 770 250 810 270
rect 770 230 780 250
rect 800 230 810 250
rect 770 210 810 230
rect 770 190 780 210
rect 800 190 810 210
rect 770 170 810 190
rect 770 150 780 170
rect 800 150 810 170
rect 770 130 810 150
rect 770 110 780 130
rect 800 110 810 130
rect 770 90 810 110
rect 770 70 780 90
rect 800 70 810 90
rect 770 50 810 70
rect 770 30 780 50
rect 800 30 810 50
rect 770 0 810 30
rect 450 -45 570 -20
rect 450 -65 460 -45
rect 480 -65 500 -45
rect 520 -65 540 -45
rect 560 -65 570 -45
rect 450 -85 570 -65
rect 365 -135 375 -115
rect 395 -135 405 -115
rect 365 -155 405 -135
rect 365 -175 375 -155
rect 395 -175 405 -155
rect 365 -195 405 -175
rect 365 -215 375 -195
rect 395 -215 405 -195
rect 365 -235 405 -215
rect 365 -255 375 -235
rect 395 -255 405 -235
rect 365 -275 405 -255
rect 365 -295 375 -275
rect 395 -295 405 -275
rect 365 -315 405 -295
rect 365 -335 375 -315
rect 395 -335 405 -315
rect 365 -355 405 -335
rect 365 -375 375 -355
rect 395 -375 405 -355
rect 365 -395 405 -375
rect 365 -415 375 -395
rect 395 -415 405 -395
rect 365 -435 405 -415
rect 365 -455 375 -435
rect 395 -455 405 -435
rect 365 -475 405 -455
rect 365 -495 375 -475
rect 395 -495 405 -475
rect 365 -505 405 -495
rect 770 -115 810 -105
rect 770 -135 780 -115
rect 800 -135 810 -115
rect 770 -155 810 -135
rect 770 -175 780 -155
rect 800 -175 810 -155
rect 770 -195 810 -175
rect 770 -215 780 -195
rect 800 -215 810 -195
rect 770 -235 810 -215
rect 770 -255 780 -235
rect 800 -255 810 -235
rect 770 -275 810 -255
rect 770 -295 780 -275
rect 800 -295 810 -275
rect 770 -315 810 -295
rect 770 -335 780 -315
rect 800 -335 810 -315
rect 770 -355 810 -335
rect 770 -375 780 -355
rect 800 -375 810 -355
rect 770 -395 810 -375
rect 770 -415 780 -395
rect 800 -415 810 -395
rect 770 -435 810 -415
rect 770 -455 780 -435
rect 800 -455 810 -435
rect 770 -475 810 -455
rect 770 -495 780 -475
rect 800 -495 810 -475
rect 770 -595 810 -495
rect -40 -635 810 -595
<< viali >>
rect -100 470 -80 490
rect 90 -65 110 -45
rect 130 -65 150 -45
rect 170 -65 190 -45
rect -100 -495 -80 -475
rect 460 -65 480 -45
rect 500 -65 520 -45
rect 540 -65 560 -45
<< metal1 >>
rect -110 490 -70 505
rect -110 470 -100 490
rect -80 470 -70 490
rect -110 455 -70 470
rect 80 -45 570 -20
rect 80 -65 90 -45
rect 110 -65 130 -45
rect 150 -65 170 -45
rect 190 -65 460 -45
rect 480 -65 500 -45
rect 520 -65 540 -45
rect 560 -65 570 -45
rect 80 -85 570 -65
rect -110 -475 -70 -460
rect -110 -495 -100 -475
rect -80 -495 -70 -475
rect -110 -510 -70 -495
<< labels >>
rlabel locali 385 -505 385 -505 5 Y
port 4 s
rlabel metal1 80 -55 80 -55 7 A
port 1 w
rlabel locali 385 630 385 630 1 VPWR
port 2 n
rlabel locali 385 -635 385 -635 5 VGND
port 3 s
rlabel metal1 -90 505 -90 505 1 VCCA
port 5 n
rlabel metal1 -90 -510 -90 -510 5 GND
port 6 s
<< end >>
