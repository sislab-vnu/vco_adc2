magic
tech sky130A
magscale 1 2
timestamp 1726562648
<< nwell >>
rect 3110 430 3190 450
rect 2030 180 2070 220
rect -690 -1760 -370 -1300
rect -680 -1810 -370 -1760
rect -690 -1860 -370 -1810
<< pwell >>
rect -930 -1780 -750 -1290
<< pdiffc >>
rect 2030 180 2070 220
<< psubdiff >>
rect -890 -1640 -790 -1620
rect -890 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -890 -1700 -790 -1680
<< nsubdiff >>
rect -570 -1640 -470 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -470 -1640
rect -570 -1700 -470 -1680
<< psubdiffcont >>
rect -860 -1680 -820 -1640
<< nsubdiffcont >>
rect -540 -1680 -500 -1640
<< locali >>
rect 180 830 990 910
rect 180 450 260 830
rect 910 450 990 830
rect 120 420 260 450
rect 120 350 180 420
rect 850 400 990 450
rect 850 350 910 400
rect 1950 350 2010 440
rect 3050 430 3190 450
rect 3050 350 3110 430
rect 3325 200 3770 350
rect -750 -980 -680 -770
rect 2190 -790 2270 80
rect 180 -890 3020 -790
rect -740 -1210 -680 -1180
rect 180 -1200 260 -890
rect -730 -1390 -690 -1210
rect 120 -1230 260 -1200
rect 120 -1300 180 -1230
rect -740 -1410 -680 -1390
rect -740 -1450 -730 -1410
rect -690 -1450 -680 -1410
rect 1140 -1450 1220 -890
rect -890 -1640 -790 -1620
rect -890 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -890 -1700 -790 -1680
rect -740 -1760 -680 -1450
rect 2060 -1460 2140 -890
rect 2940 -1200 3020 -890
rect 2880 -1240 3020 -1200
rect 2880 -1300 2940 -1240
rect -570 -1640 -470 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -470 -1640
rect -570 -1700 -470 -1680
rect 1320 -1760 1400 -1730
rect -730 -1810 -690 -1760
rect 1320 -1850 1460 -1760
rect 2320 -1840 2380 -1760
rect -740 -1940 -690 -1930
rect -730 -2060 -690 -1940
rect -740 -2190 -690 -2060
rect -740 -2220 -620 -2190
rect -740 -2280 -710 -2220
rect -650 -2280 -620 -2220
rect -740 -2310 -620 -2280
rect 360 -2360 440 -2000
rect 1320 -2360 1400 -1850
rect 360 -2460 1400 -2360
rect 2240 -1860 2380 -1840
rect 2240 -2360 2320 -1860
rect 3120 -2360 3200 -2000
rect 3670 -2360 3770 200
rect 2240 -2460 3770 -2360
rect 360 -3060 440 -2460
rect 360 -3130 590 -3060
rect 3120 -3130 3240 -3060
<< viali >>
rect 380 380 420 420
rect 3130 380 3170 420
rect 380 300 420 340
rect 3130 300 3170 340
rect 2030 180 2070 220
rect 2030 100 2070 140
rect -730 -1450 -690 -1410
rect -860 -1680 -820 -1640
rect -540 -1680 -500 -1640
rect -710 -2280 -650 -2220
<< metal1 >>
rect 360 670 3190 770
rect 360 420 440 670
rect 360 380 380 420
rect 420 380 440 420
rect 360 340 440 380
rect 360 300 380 340
rect 420 300 440 340
rect 360 280 440 300
rect 3110 420 3190 670
rect 3110 380 3130 420
rect 3170 380 3190 420
rect 3110 340 3190 380
rect 3110 300 3130 340
rect 3170 300 3190 340
rect 3110 280 3190 300
rect 2010 220 2090 240
rect 2010 210 2030 220
rect 1530 180 2030 210
rect 2070 180 2090 220
rect 1530 140 2090 180
rect 1530 110 2030 140
rect 2010 100 2030 110
rect 2070 100 2090 140
rect 2010 80 2090 100
rect -250 -680 1760 -580
rect -750 -1400 -670 -1390
rect -250 -1400 -150 -680
rect 350 -1060 450 -680
rect -750 -1410 -150 -1400
rect -750 -1450 -730 -1410
rect -690 -1450 -150 -1410
rect -750 -1460 -150 -1450
rect -750 -1470 -670 -1460
rect -890 -1640 -790 -1620
rect -890 -1680 -860 -1640
rect -820 -1680 -790 -1640
rect -890 -1700 -790 -1680
rect -570 -1640 -470 -1620
rect -570 -1680 -540 -1640
rect -500 -1680 -470 -1640
rect -570 -1700 -470 -1680
rect 1660 -1930 1760 -680
rect 1660 -2010 1960 -1930
rect -740 -2220 2850 -2190
rect -740 -2280 -710 -2220
rect -650 -2280 2850 -2220
rect -740 -2310 2850 -2280
use n_lk  n_lk_0
timestamp 1726545299
transform -1 0 1320 0 -1 -1450
box -260 -80 400 560
use n_lk  n_lk_1
timestamp 1726545299
transform -1 0 2240 0 -1 -1450
box -260 -80 400 560
use p_br1  p_br1_0
timestamp 1726477358
transform 1 0 260 0 1 80
box -260 -80 216 440
use p_br1  p_br1_1
timestamp 1726477358
transform 1 0 3190 0 1 80
box -260 -80 216 440
use p_br2  p_br2_0
timestamp 1726544869
transform 1 0 990 0 1 80
box -260 -80 580 520
use p_br2  p_br2_1
timestamp 1726544869
transform 1 0 2090 0 1 80
box -260 -80 580 520
use p_lk  p_lk_0
timestamp 1726545152
transform 1 0 260 0 1 -2010
box -260 -80 400 980
use p_lk  p_lk_1
timestamp 1726545152
transform 1 0 3020 0 1 -2010
box -260 -80 400 980
use sky130_fd_pr__res_xhigh_po_0p35_R469US  sky130_fd_pr__res_xhigh_po_0p35_R469US_0
timestamp 1726131431
transform 0 1 1848 -1 0 -3095
box -35 -1272 35 1272
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -952 -1 0 -946
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -952 -1 0 -1776
box -38 -48 314 592
<< labels >>
rlabel locali 260 910 260 910 1 VCCA
rlabel metal1 440 770 440 770 1 note_12
rlabel metal1 1700 210 1700 210 1 note_34
rlabel locali 2140 -790 2140 -790 1 add_pwr
rlabel locali 510 -3060 510 -3060 1 input_R
<< end >>
