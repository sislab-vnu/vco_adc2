* NGSPICE file created from n_lk.ext - technology: sky130A

.subckt n_lk
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5 M=2
.ends

