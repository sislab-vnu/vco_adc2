magic
tech sky130A
timestamp 1723549246
<< nwell >>
rect 30 1035 50 1055
rect 980 1035 1000 1055
rect 1460 1035 1480 1055
rect 30 995 50 1015
rect 980 995 1000 1015
rect 2005 995 2025 1015
rect 1460 955 1480 975
rect 2005 955 2025 975
rect 1450 950 1490 955
<< pwell >>
rect 20 -40 40 480
rect 8535 180 8575 260
rect 8655 220 8675 310
rect 8545 110 8565 130
rect 8545 70 8565 90
rect 7085 -625 7175 -605
rect 7085 -655 7230 -625
rect 7085 -675 7270 -655
rect 7085 -695 7175 -675
<< pdiff >>
rect 1450 950 1490 955
<< ndiffc >>
rect 8545 110 8565 130
rect 8545 70 8565 90
<< pdiffc >>
rect 30 1035 50 1055
rect 980 1035 1000 1055
rect 1460 1035 1480 1055
rect 30 995 50 1015
rect 980 995 1000 1015
rect 2005 995 2025 1015
rect 1460 955 1480 975
rect 2005 955 2025 975
<< locali >>
rect 1450 950 1490 955
rect 900 -155 940 55
rect 3765 -125 3805 55
rect 4790 -125 4830 55
rect 6630 -125 6670 55
rect 2355 -155 7050 -125
rect 7655 -155 7695 55
rect 900 -195 7695 -155
rect 2345 -225 7050 -195
rect 2345 -420 2385 -225
rect 3370 -420 3410 -225
rect 5210 -420 5250 -225
rect 6235 -420 6275 -225
<< viali >>
rect 8545 150 8565 170
rect 8545 110 8565 130
rect 8545 70 8565 90
<< metal1 >>
rect -170 785 0 835
rect 8595 785 8675 835
rect -170 -1150 -120 785
rect -70 260 0 310
rect -70 -625 -20 260
rect 20 -20 40 175
rect 8535 170 8575 260
rect 8535 150 8545 170
rect 8565 150 8575 170
rect 8535 130 8575 150
rect 8535 110 8545 130
rect 8565 110 8575 130
rect 8535 90 8575 110
rect 8535 70 8545 90
rect 8565 70 8575 90
rect 20 -70 7765 -20
rect 2275 -295 2315 -70
rect 7115 -295 7155 -70
rect 2275 -345 7155 -295
rect 8535 -625 8575 70
rect -70 -675 1445 -625
rect 7175 -675 8575 -625
rect 8625 -1150 8675 785
rect -170 -1200 1455 -1150
rect 7175 -1200 8675 -1150
use cc_inv  cc_inv_0
timestamp 1723548123
transform 1 0 60 0 1 20
box -60 -40 2805 1125
use cc_inv  cc_inv_1
timestamp 1723548123
transform 1 0 2925 0 1 20
box -60 -40 2805 1125
use cc_inv  cc_inv_2
timestamp 1723548123
transform 1 0 5790 0 1 20
box -60 -40 2805 1125
use cc_inv  cc_inv_3
timestamp 1723548123
transform -1 0 4250 0 -1 -385
box -60 -40 2805 1125
use cc_inv  cc_inv_4
timestamp 1723548123
transform -1 0 7115 0 -1 -385
box -60 -40 2805 1125
<< end >>
