magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect -580 -80 -100 440
rect 170 -80 1010 440
rect 1270 -80 2110 440
rect 2370 -90 2850 430
rect -1560 -2110 -1230 -1880
rect -510 -1930 150 -970
rect 2260 -1940 2920 -980
<< pwell >>
rect -1786 -2026 -1634 -1894
rect 464 -1054 596 -1044
rect 464 -1196 1096 -1054
rect 604 -1506 1096 -1196
rect 1374 -1364 1866 -1054
rect 1374 -1506 2006 -1364
rect 1874 -1516 2006 -1506
<< nmos >>
rect 710 -1480 810 -1080
rect 890 -1480 990 -1080
rect 1480 -1480 1580 -1080
rect 1660 -1480 1760 -1080
<< pmoshvt >>
rect -320 0 -220 360
rect 430 0 530 360
rect 610 0 710 360
rect 790 0 890 360
rect 1530 0 1630 360
rect 1710 0 1810 360
rect 1890 0 1990 360
rect 2630 -10 2730 350
rect -250 -1850 -150 -1050
rect -70 -1850 30 -1050
rect 2520 -1860 2620 -1060
rect 2700 -1860 2800 -1060
<< ndiff >>
rect 630 -1113 710 -1080
rect 630 -1147 653 -1113
rect 687 -1147 710 -1113
rect 630 -1193 710 -1147
rect 630 -1227 653 -1193
rect 687 -1227 710 -1193
rect 630 -1273 710 -1227
rect 630 -1307 653 -1273
rect 687 -1307 710 -1273
rect 630 -1353 710 -1307
rect 630 -1387 653 -1353
rect 687 -1387 710 -1353
rect 630 -1480 710 -1387
rect 810 -1113 890 -1080
rect 810 -1147 833 -1113
rect 867 -1147 890 -1113
rect 810 -1193 890 -1147
rect 810 -1227 833 -1193
rect 867 -1227 890 -1193
rect 810 -1273 890 -1227
rect 810 -1307 833 -1273
rect 867 -1307 890 -1273
rect 810 -1353 890 -1307
rect 810 -1387 833 -1353
rect 867 -1387 890 -1353
rect 810 -1480 890 -1387
rect 990 -1113 1070 -1080
rect 990 -1147 1013 -1113
rect 1047 -1147 1070 -1113
rect 990 -1193 1070 -1147
rect 990 -1227 1013 -1193
rect 1047 -1227 1070 -1193
rect 990 -1273 1070 -1227
rect 990 -1307 1013 -1273
rect 1047 -1307 1070 -1273
rect 990 -1353 1070 -1307
rect 990 -1387 1013 -1353
rect 1047 -1387 1070 -1353
rect 990 -1480 1070 -1387
rect 1400 -1173 1480 -1080
rect 1400 -1207 1423 -1173
rect 1457 -1207 1480 -1173
rect 1400 -1253 1480 -1207
rect 1400 -1287 1423 -1253
rect 1457 -1287 1480 -1253
rect 1400 -1333 1480 -1287
rect 1400 -1367 1423 -1333
rect 1457 -1367 1480 -1333
rect 1400 -1413 1480 -1367
rect 1400 -1447 1423 -1413
rect 1457 -1447 1480 -1413
rect 1400 -1480 1480 -1447
rect 1580 -1173 1660 -1080
rect 1580 -1207 1603 -1173
rect 1637 -1207 1660 -1173
rect 1580 -1253 1660 -1207
rect 1580 -1287 1603 -1253
rect 1637 -1287 1660 -1253
rect 1580 -1333 1660 -1287
rect 1580 -1367 1603 -1333
rect 1637 -1367 1660 -1333
rect 1580 -1413 1660 -1367
rect 1580 -1447 1603 -1413
rect 1637 -1447 1660 -1413
rect 1580 -1480 1660 -1447
rect 1760 -1173 1840 -1080
rect 1760 -1207 1783 -1173
rect 1817 -1207 1840 -1173
rect 1760 -1253 1840 -1207
rect 1760 -1287 1783 -1253
rect 1817 -1287 1840 -1253
rect 1760 -1333 1840 -1287
rect 1760 -1367 1783 -1333
rect 1817 -1367 1840 -1333
rect 1760 -1413 1840 -1367
rect 1760 -1447 1783 -1413
rect 1817 -1447 1840 -1413
rect 1760 -1480 1840 -1447
<< pdiff >>
rect -400 337 -320 360
rect -400 303 -377 337
rect -343 303 -320 337
rect -400 257 -320 303
rect -400 223 -377 257
rect -343 223 -320 257
rect -400 177 -320 223
rect -400 143 -377 177
rect -343 143 -320 177
rect -400 97 -320 143
rect -400 63 -377 97
rect -343 63 -320 97
rect -400 0 -320 63
rect -220 337 -140 360
rect -220 303 -197 337
rect -163 303 -140 337
rect -220 257 -140 303
rect 350 337 430 360
rect 350 303 373 337
rect 407 303 430 337
rect -220 223 -197 257
rect -163 223 -140 257
rect -220 177 -140 223
rect -220 143 -197 177
rect -163 143 -140 177
rect -220 97 -140 143
rect -220 63 -197 97
rect -163 63 -140 97
rect -220 0 -140 63
rect 350 257 430 303
rect 350 223 373 257
rect 407 223 430 257
rect 350 177 430 223
rect 350 143 373 177
rect 407 143 430 177
rect 350 97 430 143
rect 350 63 373 97
rect 407 63 430 97
rect 350 0 430 63
rect 530 337 610 360
rect 530 303 553 337
rect 587 303 610 337
rect 530 257 610 303
rect 530 223 553 257
rect 587 223 610 257
rect 530 177 610 223
rect 530 143 553 177
rect 587 143 610 177
rect 530 97 610 143
rect 530 63 553 97
rect 587 63 610 97
rect 530 0 610 63
rect 710 337 790 360
rect 710 303 733 337
rect 767 303 790 337
rect 710 257 790 303
rect 710 223 733 257
rect 767 223 790 257
rect 710 177 790 223
rect 710 143 733 177
rect 767 143 790 177
rect 710 97 790 143
rect 710 63 733 97
rect 767 63 790 97
rect 710 0 790 63
rect 890 337 970 360
rect 890 303 913 337
rect 947 303 970 337
rect 890 257 970 303
rect 1450 337 1530 360
rect 1450 303 1473 337
rect 1507 303 1530 337
rect 890 223 913 257
rect 947 223 970 257
rect 890 177 970 223
rect 890 143 913 177
rect 947 143 970 177
rect 890 97 970 143
rect 890 63 913 97
rect 947 63 970 97
rect 890 0 970 63
rect 1450 257 1530 303
rect 1450 223 1473 257
rect 1507 223 1530 257
rect 1450 177 1530 223
rect 1450 143 1473 177
rect 1507 143 1530 177
rect 1450 97 1530 143
rect 1450 63 1473 97
rect 1507 63 1530 97
rect 1450 0 1530 63
rect 1630 337 1710 360
rect 1630 303 1653 337
rect 1687 303 1710 337
rect 1630 257 1710 303
rect 1630 223 1653 257
rect 1687 223 1710 257
rect 1630 177 1710 223
rect 1630 143 1653 177
rect 1687 143 1710 177
rect 1630 97 1710 143
rect 1630 63 1653 97
rect 1687 63 1710 97
rect 1630 0 1710 63
rect 1810 337 1890 360
rect 1810 303 1833 337
rect 1867 303 1890 337
rect 1810 257 1890 303
rect 1810 223 1833 257
rect 1867 223 1890 257
rect 1810 177 1890 223
rect 1810 143 1833 177
rect 1867 143 1890 177
rect 1810 97 1890 143
rect 1810 63 1833 97
rect 1867 63 1890 97
rect 1810 0 1890 63
rect 1990 337 2070 360
rect 1990 303 2013 337
rect 2047 303 2070 337
rect 1990 257 2070 303
rect 2550 327 2630 350
rect 2550 293 2573 327
rect 2607 293 2630 327
rect 1990 223 2013 257
rect 2047 223 2070 257
rect 1990 177 2070 223
rect 1990 143 2013 177
rect 2047 143 2070 177
rect 1990 97 2070 143
rect 1990 63 2013 97
rect 2047 63 2070 97
rect 1990 0 2070 63
rect 2550 247 2630 293
rect 2550 213 2573 247
rect 2607 213 2630 247
rect 2550 167 2630 213
rect 2550 133 2573 167
rect 2607 133 2630 167
rect 2550 87 2630 133
rect 2550 53 2573 87
rect 2607 53 2630 87
rect 2550 -10 2630 53
rect 2730 327 2810 350
rect 2730 293 2753 327
rect 2787 293 2810 327
rect 2730 247 2810 293
rect 2730 213 2753 247
rect 2787 213 2810 247
rect 2730 167 2810 213
rect 2730 133 2753 167
rect 2787 133 2810 167
rect 2730 87 2810 133
rect 2730 53 2753 87
rect 2787 53 2810 87
rect 2730 -10 2810 53
rect -330 -1073 -250 -1050
rect -330 -1107 -307 -1073
rect -273 -1107 -250 -1073
rect -330 -1153 -250 -1107
rect -330 -1187 -307 -1153
rect -273 -1187 -250 -1153
rect -330 -1233 -250 -1187
rect -330 -1267 -307 -1233
rect -273 -1267 -250 -1233
rect -330 -1313 -250 -1267
rect -330 -1347 -307 -1313
rect -273 -1347 -250 -1313
rect -330 -1393 -250 -1347
rect -330 -1427 -307 -1393
rect -273 -1427 -250 -1393
rect -330 -1473 -250 -1427
rect -330 -1507 -307 -1473
rect -273 -1507 -250 -1473
rect -330 -1553 -250 -1507
rect -330 -1587 -307 -1553
rect -273 -1587 -250 -1553
rect -330 -1633 -250 -1587
rect -330 -1667 -307 -1633
rect -273 -1667 -250 -1633
rect -330 -1713 -250 -1667
rect -330 -1747 -307 -1713
rect -273 -1747 -250 -1713
rect -330 -1793 -250 -1747
rect -330 -1827 -307 -1793
rect -273 -1827 -250 -1793
rect -330 -1850 -250 -1827
rect -150 -1073 -70 -1050
rect -150 -1107 -127 -1073
rect -93 -1107 -70 -1073
rect -150 -1153 -70 -1107
rect -150 -1187 -127 -1153
rect -93 -1187 -70 -1153
rect -150 -1233 -70 -1187
rect -150 -1267 -127 -1233
rect -93 -1267 -70 -1233
rect -150 -1313 -70 -1267
rect -150 -1347 -127 -1313
rect -93 -1347 -70 -1313
rect -150 -1393 -70 -1347
rect -150 -1427 -127 -1393
rect -93 -1427 -70 -1393
rect -150 -1473 -70 -1427
rect -150 -1507 -127 -1473
rect -93 -1507 -70 -1473
rect -150 -1553 -70 -1507
rect -150 -1587 -127 -1553
rect -93 -1587 -70 -1553
rect -150 -1633 -70 -1587
rect -150 -1667 -127 -1633
rect -93 -1667 -70 -1633
rect -150 -1713 -70 -1667
rect -150 -1747 -127 -1713
rect -93 -1747 -70 -1713
rect -150 -1793 -70 -1747
rect -150 -1827 -127 -1793
rect -93 -1827 -70 -1793
rect -150 -1850 -70 -1827
rect 30 -1073 110 -1050
rect 30 -1107 53 -1073
rect 87 -1107 110 -1073
rect 30 -1153 110 -1107
rect 30 -1187 53 -1153
rect 87 -1187 110 -1153
rect 30 -1233 110 -1187
rect 30 -1267 53 -1233
rect 87 -1267 110 -1233
rect 30 -1313 110 -1267
rect 30 -1347 53 -1313
rect 87 -1347 110 -1313
rect 30 -1393 110 -1347
rect 30 -1427 53 -1393
rect 87 -1427 110 -1393
rect 30 -1473 110 -1427
rect 30 -1507 53 -1473
rect 87 -1507 110 -1473
rect 2440 -1083 2520 -1060
rect 2440 -1117 2463 -1083
rect 2497 -1117 2520 -1083
rect 2440 -1163 2520 -1117
rect 2440 -1197 2463 -1163
rect 2497 -1197 2520 -1163
rect 2440 -1243 2520 -1197
rect 2440 -1277 2463 -1243
rect 2497 -1277 2520 -1243
rect 2440 -1323 2520 -1277
rect 2440 -1357 2463 -1323
rect 2497 -1357 2520 -1323
rect 30 -1553 110 -1507
rect 30 -1587 53 -1553
rect 87 -1587 110 -1553
rect 30 -1633 110 -1587
rect 30 -1667 53 -1633
rect 87 -1667 110 -1633
rect 2440 -1403 2520 -1357
rect 2440 -1437 2463 -1403
rect 2497 -1437 2520 -1403
rect 2440 -1483 2520 -1437
rect 2440 -1517 2463 -1483
rect 2497 -1517 2520 -1483
rect 2440 -1563 2520 -1517
rect 2440 -1597 2463 -1563
rect 2497 -1597 2520 -1563
rect 2440 -1643 2520 -1597
rect 30 -1713 110 -1667
rect 30 -1747 53 -1713
rect 87 -1747 110 -1713
rect 30 -1793 110 -1747
rect 30 -1827 53 -1793
rect 87 -1827 110 -1793
rect 30 -1850 110 -1827
rect 2440 -1677 2463 -1643
rect 2497 -1677 2520 -1643
rect 2440 -1723 2520 -1677
rect 2440 -1757 2463 -1723
rect 2497 -1757 2520 -1723
rect 2440 -1803 2520 -1757
rect 2440 -1837 2463 -1803
rect 2497 -1837 2520 -1803
rect 2440 -1860 2520 -1837
rect 2620 -1083 2700 -1060
rect 2620 -1117 2643 -1083
rect 2677 -1117 2700 -1083
rect 2620 -1163 2700 -1117
rect 2620 -1197 2643 -1163
rect 2677 -1197 2700 -1163
rect 2620 -1243 2700 -1197
rect 2620 -1277 2643 -1243
rect 2677 -1277 2700 -1243
rect 2620 -1323 2700 -1277
rect 2620 -1357 2643 -1323
rect 2677 -1357 2700 -1323
rect 2620 -1403 2700 -1357
rect 2620 -1437 2643 -1403
rect 2677 -1437 2700 -1403
rect 2620 -1483 2700 -1437
rect 2620 -1517 2643 -1483
rect 2677 -1517 2700 -1483
rect 2620 -1563 2700 -1517
rect 2620 -1597 2643 -1563
rect 2677 -1597 2700 -1563
rect 2620 -1643 2700 -1597
rect 2620 -1677 2643 -1643
rect 2677 -1677 2700 -1643
rect 2620 -1723 2700 -1677
rect 2620 -1757 2643 -1723
rect 2677 -1757 2700 -1723
rect 2620 -1803 2700 -1757
rect 2620 -1837 2643 -1803
rect 2677 -1837 2700 -1803
rect 2620 -1860 2700 -1837
rect 2800 -1083 2880 -1060
rect 2800 -1117 2823 -1083
rect 2857 -1117 2880 -1083
rect 2800 -1163 2880 -1117
rect 2800 -1197 2823 -1163
rect 2857 -1197 2880 -1163
rect 2800 -1243 2880 -1197
rect 2800 -1277 2823 -1243
rect 2857 -1277 2880 -1243
rect 2800 -1323 2880 -1277
rect 2800 -1357 2823 -1323
rect 2857 -1357 2880 -1323
rect 2800 -1403 2880 -1357
rect 2800 -1437 2823 -1403
rect 2857 -1437 2880 -1403
rect 2800 -1483 2880 -1437
rect 2800 -1517 2823 -1483
rect 2857 -1517 2880 -1483
rect 2800 -1563 2880 -1517
rect 2800 -1597 2823 -1563
rect 2857 -1597 2880 -1563
rect 2800 -1643 2880 -1597
rect 2800 -1677 2823 -1643
rect 2857 -1677 2880 -1643
rect 2800 -1723 2880 -1677
rect 2800 -1757 2823 -1723
rect 2857 -1757 2880 -1723
rect 2800 -1803 2880 -1757
rect 2800 -1837 2823 -1803
rect 2857 -1837 2880 -1803
rect 2800 -1860 2880 -1837
<< ndiffc >>
rect 653 -1147 687 -1113
rect 653 -1227 687 -1193
rect 653 -1307 687 -1273
rect 653 -1387 687 -1353
rect 833 -1147 867 -1113
rect 833 -1227 867 -1193
rect 833 -1307 867 -1273
rect 833 -1387 867 -1353
rect 1013 -1147 1047 -1113
rect 1013 -1227 1047 -1193
rect 1013 -1307 1047 -1273
rect 1013 -1387 1047 -1353
rect 1423 -1207 1457 -1173
rect 1423 -1287 1457 -1253
rect 1423 -1367 1457 -1333
rect 1423 -1447 1457 -1413
rect 1603 -1207 1637 -1173
rect 1603 -1287 1637 -1253
rect 1603 -1367 1637 -1333
rect 1603 -1447 1637 -1413
rect 1783 -1207 1817 -1173
rect 1783 -1287 1817 -1253
rect 1783 -1367 1817 -1333
rect 1783 -1447 1817 -1413
<< pdiffc >>
rect -377 303 -343 337
rect -377 223 -343 257
rect -377 143 -343 177
rect -377 63 -343 97
rect -197 303 -163 337
rect 373 303 407 337
rect -197 223 -163 257
rect -197 143 -163 177
rect -197 63 -163 97
rect 373 223 407 257
rect 373 143 407 177
rect 373 63 407 97
rect 553 303 587 337
rect 553 223 587 257
rect 553 143 587 177
rect 553 63 587 97
rect 733 303 767 337
rect 733 223 767 257
rect 733 143 767 177
rect 733 63 767 97
rect 913 303 947 337
rect 1473 303 1507 337
rect 913 223 947 257
rect 913 143 947 177
rect 913 63 947 97
rect 1473 223 1507 257
rect 1473 143 1507 177
rect 1473 63 1507 97
rect 1653 303 1687 337
rect 1653 223 1687 257
rect 1653 143 1687 177
rect 1653 63 1687 97
rect 1833 303 1867 337
rect 1833 223 1867 257
rect 1833 143 1867 177
rect 1833 63 1867 97
rect 2013 303 2047 337
rect 2573 293 2607 327
rect 2013 223 2047 257
rect 2013 143 2047 177
rect 2013 63 2047 97
rect 2573 213 2607 247
rect 2573 133 2607 167
rect 2573 53 2607 87
rect 2753 293 2787 327
rect 2753 213 2787 247
rect 2753 133 2787 167
rect 2753 53 2787 87
rect -307 -1107 -273 -1073
rect -307 -1187 -273 -1153
rect -307 -1267 -273 -1233
rect -307 -1347 -273 -1313
rect -307 -1427 -273 -1393
rect -307 -1507 -273 -1473
rect -307 -1587 -273 -1553
rect -307 -1667 -273 -1633
rect -307 -1747 -273 -1713
rect -307 -1827 -273 -1793
rect -127 -1107 -93 -1073
rect -127 -1187 -93 -1153
rect -127 -1267 -93 -1233
rect -127 -1347 -93 -1313
rect -127 -1427 -93 -1393
rect -127 -1507 -93 -1473
rect -127 -1587 -93 -1553
rect -127 -1667 -93 -1633
rect -127 -1747 -93 -1713
rect -127 -1827 -93 -1793
rect 53 -1107 87 -1073
rect 53 -1187 87 -1153
rect 53 -1267 87 -1233
rect 53 -1347 87 -1313
rect 53 -1427 87 -1393
rect 53 -1507 87 -1473
rect 2463 -1117 2497 -1083
rect 2463 -1197 2497 -1163
rect 2463 -1277 2497 -1243
rect 2463 -1357 2497 -1323
rect 53 -1587 87 -1553
rect 53 -1667 87 -1633
rect 2463 -1437 2497 -1403
rect 2463 -1517 2497 -1483
rect 2463 -1597 2497 -1563
rect 53 -1747 87 -1713
rect 53 -1827 87 -1793
rect 2463 -1677 2497 -1643
rect 2463 -1757 2497 -1723
rect 2463 -1837 2497 -1803
rect 2643 -1117 2677 -1083
rect 2643 -1197 2677 -1163
rect 2643 -1277 2677 -1243
rect 2643 -1357 2677 -1323
rect 2643 -1437 2677 -1403
rect 2643 -1517 2677 -1483
rect 2643 -1597 2677 -1563
rect 2643 -1677 2677 -1643
rect 2643 -1757 2677 -1723
rect 2643 -1837 2677 -1803
rect 2823 -1117 2857 -1083
rect 2823 -1197 2857 -1163
rect 2823 -1277 2857 -1243
rect 2823 -1357 2857 -1323
rect 2823 -1437 2857 -1403
rect 2823 -1517 2857 -1483
rect 2823 -1597 2857 -1563
rect 2823 -1677 2857 -1643
rect 2823 -1757 2857 -1723
rect 2823 -1837 2857 -1803
<< psubdiff >>
rect 490 -1103 570 -1070
rect 490 -1137 513 -1103
rect 547 -1137 570 -1103
rect 490 -1170 570 -1137
rect 1900 -1423 1980 -1390
rect 1900 -1457 1923 -1423
rect 1957 -1457 1980 -1423
rect 1900 -1490 1980 -1457
rect -1760 -1943 -1660 -1920
rect -1760 -1977 -1727 -1943
rect -1693 -1977 -1660 -1943
rect -1760 -2000 -1660 -1977
<< nsubdiff >>
rect -540 327 -460 360
rect -540 293 -517 327
rect -483 293 -460 327
rect -540 260 -460 293
rect 210 337 290 370
rect 210 303 233 337
rect 267 303 290 337
rect 210 270 290 303
rect 1310 337 1390 370
rect 1310 303 1333 337
rect 1367 303 1390 337
rect 1310 270 1390 303
rect 2410 327 2490 360
rect 2410 293 2433 327
rect 2467 293 2490 327
rect 2410 260 2490 293
rect -470 -1073 -390 -1040
rect -470 -1107 -447 -1073
rect -413 -1107 -390 -1073
rect -470 -1140 -390 -1107
rect 2300 -1103 2380 -1070
rect 2300 -1137 2323 -1103
rect 2357 -1137 2380 -1103
rect 2300 -1170 2380 -1137
rect -1480 -1923 -1380 -1900
rect -1480 -1957 -1447 -1923
rect -1413 -1957 -1380 -1923
rect -1480 -1980 -1380 -1957
<< psubdiffcont >>
rect 513 -1137 547 -1103
rect 1923 -1457 1957 -1423
rect -1727 -1977 -1693 -1943
<< nsubdiffcont >>
rect -517 293 -483 327
rect 233 303 267 337
rect 1333 303 1367 337
rect 2433 293 2467 327
rect -447 -1107 -413 -1073
rect 2323 -1137 2357 -1103
rect -1447 -1957 -1413 -1923
<< poly >>
rect -320 507 -220 540
rect -320 473 -267 507
rect -233 473 -220 507
rect -320 360 -220 473
rect 430 507 890 540
rect 430 473 503 507
rect 537 473 603 507
rect 637 473 890 507
rect 430 440 890 473
rect 430 360 530 440
rect 610 360 710 440
rect 790 360 890 440
rect 1530 507 1990 540
rect 1530 473 1563 507
rect 1597 473 1743 507
rect 1777 473 1923 507
rect 1957 473 1990 507
rect 1530 440 1990 473
rect 1530 360 1630 440
rect 1710 360 1810 440
rect 1890 360 1990 440
rect 2630 497 2730 530
rect 2630 463 2663 497
rect 2697 463 2730 497
rect 2630 350 2730 463
rect -320 -80 -220 0
rect 430 -80 530 0
rect 610 -80 710 0
rect 790 -80 890 0
rect 1530 -80 1630 0
rect 1710 -80 1810 0
rect 1890 -80 1990 0
rect 2630 -90 2730 -10
rect -250 -1050 -150 -970
rect -70 -1050 30 -970
rect 710 -1080 810 -1000
rect 890 -1080 990 -1000
rect 1480 -1080 1580 -1000
rect 1660 -1080 1760 -1000
rect 2520 -1060 2620 -980
rect 2700 -1060 2800 -980
rect 710 -1560 810 -1480
rect 890 -1560 990 -1480
rect 710 -1593 990 -1560
rect 710 -1627 783 -1593
rect 817 -1627 883 -1593
rect 917 -1627 990 -1593
rect 710 -1660 990 -1627
rect 1480 -1560 1580 -1480
rect 1660 -1560 1760 -1480
rect 1480 -1593 1760 -1560
rect 1480 -1627 1563 -1593
rect 1597 -1627 1653 -1593
rect 1687 -1627 1760 -1593
rect 1480 -1660 1760 -1627
rect -250 -1930 -150 -1850
rect -70 -1930 30 -1850
rect -250 -1963 30 -1930
rect -250 -1997 -237 -1963
rect -203 -1997 -17 -1963
rect 17 -1997 30 -1963
rect -250 -2030 30 -1997
rect 2520 -1940 2620 -1860
rect 2700 -1940 2800 -1860
rect 2520 -1973 2800 -1940
rect 2520 -2007 2533 -1973
rect 2567 -2007 2753 -1973
rect 2787 -2007 2800 -1973
rect 2520 -2040 2800 -2007
<< polycont >>
rect -267 473 -233 507
rect 503 473 537 507
rect 603 473 637 507
rect 1563 473 1597 507
rect 1743 473 1777 507
rect 1923 473 1957 507
rect 2663 463 2697 497
rect 783 -1627 817 -1593
rect 883 -1627 917 -1593
rect 1563 -1627 1597 -1593
rect 1653 -1627 1687 -1593
rect -237 -1997 -203 -1963
rect -17 -1997 17 -1963
rect 2533 -2007 2567 -1973
rect 2753 -2007 2787 -1973
<< locali >>
rect -540 660 790 740
rect -540 327 -460 660
rect -540 293 -517 327
rect -483 293 -460 327
rect -540 260 -460 293
rect -400 337 -320 660
rect -280 507 -220 540
rect -280 473 -267 507
rect -233 473 -220 507
rect -280 440 -220 473
rect -400 303 -377 337
rect -343 303 -320 337
rect -400 257 -320 303
rect -400 223 -377 257
rect -343 223 -320 257
rect -400 177 -320 223
rect -400 143 -377 177
rect -343 143 -320 177
rect -400 97 -320 143
rect -400 63 -377 97
rect -343 63 -320 97
rect -400 0 -320 63
rect -220 337 -140 360
rect -220 303 -197 337
rect -163 303 -140 337
rect -220 257 -140 303
rect 210 337 290 660
rect 470 507 670 540
rect 470 473 503 507
rect 537 473 603 507
rect 637 473 670 507
rect 470 440 670 473
rect 210 303 233 337
rect 267 303 290 337
rect 210 270 290 303
rect 350 337 430 360
rect 350 303 373 337
rect 407 303 430 337
rect -220 223 -197 257
rect -163 223 -140 257
rect -220 177 -140 223
rect -220 143 -197 177
rect -163 143 -140 177
rect -220 97 -140 143
rect -220 63 -197 97
rect -163 63 -140 97
rect -220 0 -140 63
rect 350 257 430 303
rect 350 223 373 257
rect 407 223 430 257
rect 350 177 430 223
rect 350 143 373 177
rect 407 143 430 177
rect 350 97 430 143
rect 350 63 373 97
rect 407 63 430 97
rect 350 0 430 63
rect 530 337 610 360
rect 530 303 553 337
rect 587 303 610 337
rect 530 257 610 303
rect 530 223 553 257
rect 587 223 610 257
rect 530 177 610 223
rect 530 143 553 177
rect 587 143 610 177
rect 530 97 610 143
rect 530 63 553 97
rect 587 63 610 97
rect 530 0 610 63
rect 710 337 790 660
rect 1530 507 1990 540
rect 1530 473 1563 507
rect 1597 473 1743 507
rect 1777 473 1923 507
rect 1957 473 1990 507
rect 1530 440 1990 473
rect 2630 497 2730 530
rect 2630 463 2663 497
rect 2697 463 2730 497
rect 2630 430 2730 463
rect 710 303 733 337
rect 767 303 790 337
rect 710 257 790 303
rect 710 223 733 257
rect 767 223 790 257
rect 710 177 790 223
rect 710 143 733 177
rect 767 143 790 177
rect 710 97 790 143
rect 710 63 733 97
rect 767 63 790 97
rect 710 0 790 63
rect 890 337 970 360
rect 890 303 913 337
rect 947 303 970 337
rect 890 257 970 303
rect 890 223 913 257
rect 947 223 970 257
rect 890 177 970 223
rect 890 143 913 177
rect 947 143 970 177
rect 890 97 970 143
rect 890 63 913 97
rect 947 63 970 97
rect 890 -150 970 63
rect 1310 337 1390 370
rect 1310 303 1333 337
rect 1367 303 1390 337
rect 1310 -150 1390 303
rect 1450 337 1530 360
rect 1450 303 1473 337
rect 1507 303 1530 337
rect 1450 257 1530 303
rect 1450 223 1473 257
rect 1507 223 1530 257
rect 1450 177 1530 223
rect 1450 143 1473 177
rect 1507 143 1530 177
rect 1450 97 1530 143
rect 1450 63 1473 97
rect 1507 63 1530 97
rect 1450 -150 1530 63
rect 890 -230 1530 -150
rect 1630 337 1710 360
rect 1630 303 1653 337
rect 1687 303 1710 337
rect 1630 257 1710 303
rect 1630 223 1653 257
rect 1687 223 1710 257
rect 1630 177 1710 223
rect 1630 143 1653 177
rect 1687 143 1710 177
rect 1630 97 1710 143
rect 1630 63 1653 97
rect 1687 63 1710 97
rect 1630 -540 1710 63
rect 1810 337 1890 360
rect 1810 303 1833 337
rect 1867 303 1890 337
rect 1810 257 1890 303
rect 1810 223 1833 257
rect 1867 223 1890 257
rect 1810 177 1890 223
rect 1810 143 1833 177
rect 1867 143 1890 177
rect 1810 97 1890 143
rect 1810 63 1833 97
rect 1867 63 1890 97
rect 1810 0 1890 63
rect 1990 337 2070 360
rect 1990 303 2013 337
rect 2047 303 2070 337
rect 1990 257 2070 303
rect 2410 327 2490 360
rect 2410 293 2433 327
rect 2467 293 2490 327
rect 2410 260 2490 293
rect 2550 327 2630 350
rect 2550 293 2573 327
rect 2607 293 2630 327
rect 1990 223 2013 257
rect 2047 223 2070 257
rect 1990 177 2070 223
rect 1990 143 2013 177
rect 2047 143 2070 177
rect 1990 97 2070 143
rect 1990 63 2013 97
rect 2047 63 2070 97
rect 1990 0 2070 63
rect 2550 247 2630 293
rect 2550 213 2573 247
rect 2607 213 2630 247
rect 2550 167 2630 213
rect 2550 133 2573 167
rect 2607 133 2630 167
rect 2550 87 2630 133
rect 2550 53 2573 87
rect 2607 53 2630 87
rect 2550 -10 2630 53
rect 2730 327 2810 350
rect 2730 293 2753 327
rect 2787 293 2810 327
rect 2730 247 2810 293
rect 2730 213 2753 247
rect 2787 213 2810 247
rect 2730 167 2810 213
rect 2730 133 2753 167
rect 2787 133 2810 167
rect 2730 90 2810 133
rect 2730 87 3220 90
rect 2730 53 2753 87
rect 2787 53 3220 87
rect 2730 -10 3220 53
rect 10 -640 2380 -540
rect 10 -740 110 -640
rect -470 -840 110 -740
rect -470 -1073 -390 -840
rect -470 -1107 -447 -1073
rect -413 -1107 -390 -1073
rect -470 -1140 -390 -1107
rect -330 -1073 -250 -1050
rect -330 -1107 -307 -1073
rect -273 -1107 -250 -1073
rect -330 -1153 -250 -1107
rect -330 -1187 -307 -1153
rect -273 -1187 -250 -1153
rect -330 -1233 -250 -1187
rect -330 -1267 -307 -1233
rect -273 -1267 -250 -1233
rect -330 -1313 -250 -1267
rect -330 -1347 -307 -1313
rect -273 -1347 -250 -1313
rect -330 -1393 -250 -1347
rect -330 -1427 -307 -1393
rect -273 -1427 -250 -1393
rect -330 -1473 -250 -1427
rect -330 -1507 -307 -1473
rect -273 -1507 -250 -1473
rect -1600 -1523 -1560 -1520
rect -1600 -1557 -1597 -1523
rect -1563 -1557 -1560 -1523
rect -1600 -1560 -1560 -1557
rect -330 -1553 -250 -1507
rect -330 -1587 -307 -1553
rect -273 -1587 -250 -1553
rect -330 -1633 -250 -1587
rect -330 -1667 -307 -1633
rect -273 -1667 -250 -1633
rect -330 -1713 -250 -1667
rect -1760 -1943 -1660 -1920
rect -1760 -1977 -1727 -1943
rect -1693 -1977 -1660 -1943
rect -1760 -2000 -1660 -1977
rect -1590 -2020 -1550 -1720
rect -330 -1747 -307 -1713
rect -273 -1747 -250 -1713
rect -330 -1793 -250 -1747
rect -330 -1827 -307 -1793
rect -273 -1827 -250 -1793
rect -330 -1850 -250 -1827
rect -150 -1073 -70 -1050
rect -150 -1107 -127 -1073
rect -93 -1107 -70 -1073
rect -150 -1153 -70 -1107
rect -150 -1187 -127 -1153
rect -93 -1187 -70 -1153
rect -150 -1233 -70 -1187
rect -150 -1267 -127 -1233
rect -93 -1267 -70 -1233
rect -150 -1313 -70 -1267
rect -150 -1347 -127 -1313
rect -93 -1347 -70 -1313
rect -150 -1393 -70 -1347
rect -150 -1427 -127 -1393
rect -93 -1427 -70 -1393
rect -150 -1473 -70 -1427
rect -150 -1507 -127 -1473
rect -93 -1507 -70 -1473
rect -150 -1553 -70 -1507
rect -150 -1587 -127 -1553
rect -93 -1587 -70 -1553
rect -150 -1633 -70 -1587
rect -150 -1667 -127 -1633
rect -93 -1667 -70 -1633
rect -150 -1713 -70 -1667
rect -150 -1747 -127 -1713
rect -93 -1747 -70 -1713
rect -150 -1793 -70 -1747
rect -150 -1827 -127 -1793
rect -93 -1827 -70 -1793
rect -1480 -1923 -1380 -1900
rect -1480 -1957 -1447 -1923
rect -1413 -1957 -1380 -1923
rect -250 -1940 -190 -1930
rect -1480 -1980 -1380 -1957
rect -1110 -1963 -190 -1940
rect -1110 -1997 -237 -1963
rect -203 -1997 -190 -1963
rect -1110 -2020 -190 -1997
rect -1590 -2100 -1030 -2020
rect -250 -2030 -190 -2020
rect -1590 -2180 -1550 -2100
rect -150 -2170 -70 -1827
rect 30 -1073 110 -840
rect 30 -1107 53 -1073
rect 87 -1107 110 -1073
rect 30 -1153 110 -1107
rect 30 -1187 53 -1153
rect 87 -1187 110 -1153
rect 490 -1103 570 -1070
rect 490 -1137 513 -1103
rect 547 -1137 570 -1103
rect 490 -1170 570 -1137
rect 630 -1113 710 -1080
rect 630 -1147 653 -1113
rect 687 -1147 710 -1113
rect 30 -1233 110 -1187
rect 30 -1267 53 -1233
rect 87 -1267 110 -1233
rect 30 -1313 110 -1267
rect 30 -1347 53 -1313
rect 87 -1347 110 -1313
rect 30 -1393 110 -1347
rect 30 -1427 53 -1393
rect 87 -1427 110 -1393
rect 30 -1473 110 -1427
rect 30 -1507 53 -1473
rect 87 -1507 110 -1473
rect 30 -1553 110 -1507
rect 30 -1587 53 -1553
rect 87 -1587 110 -1553
rect 30 -1633 110 -1587
rect 30 -1667 53 -1633
rect 87 -1667 110 -1633
rect 30 -1713 110 -1667
rect 30 -1747 53 -1713
rect 87 -1747 110 -1713
rect 30 -1793 110 -1747
rect 30 -1827 53 -1793
rect 87 -1827 110 -1793
rect 30 -1850 110 -1827
rect 630 -1193 710 -1147
rect 630 -1227 653 -1193
rect 687 -1227 710 -1193
rect 630 -1273 710 -1227
rect 630 -1307 653 -1273
rect 687 -1307 710 -1273
rect 630 -1353 710 -1307
rect 630 -1387 653 -1353
rect 687 -1387 710 -1353
rect -30 -1963 30 -1930
rect -30 -1997 -17 -1963
rect 17 -1997 30 -1963
rect -30 -2030 30 -1997
rect 630 -2170 710 -1387
rect 810 -1113 890 -640
rect 810 -1147 833 -1113
rect 867 -1147 890 -1113
rect 810 -1193 890 -1147
rect 810 -1227 833 -1193
rect 867 -1227 890 -1193
rect 810 -1273 890 -1227
rect 810 -1307 833 -1273
rect 867 -1307 890 -1273
rect 810 -1353 890 -1307
rect 810 -1387 833 -1353
rect 867 -1387 890 -1353
rect 810 -1480 890 -1387
rect 990 -1113 1070 -1080
rect 990 -1147 1013 -1113
rect 1047 -1147 1070 -1113
rect 990 -1193 1070 -1147
rect 990 -1227 1013 -1193
rect 1047 -1227 1070 -1193
rect 990 -1273 1070 -1227
rect 990 -1307 1013 -1273
rect 1047 -1307 1070 -1273
rect 990 -1353 1070 -1307
rect 990 -1387 1013 -1353
rect 1047 -1387 1070 -1353
rect 990 -1480 1070 -1387
rect 1400 -1173 1480 -1080
rect 1400 -1207 1423 -1173
rect 1457 -1207 1480 -1173
rect 1400 -1253 1480 -1207
rect 1400 -1287 1423 -1253
rect 1457 -1287 1480 -1253
rect 1400 -1333 1480 -1287
rect 1400 -1367 1423 -1333
rect 1457 -1367 1480 -1333
rect 1400 -1413 1480 -1367
rect 1400 -1447 1423 -1413
rect 1457 -1447 1480 -1413
rect 1400 -1480 1480 -1447
rect 1580 -1173 1660 -640
rect 2300 -740 2380 -640
rect 2300 -840 2520 -740
rect 1580 -1207 1603 -1173
rect 1637 -1207 1660 -1173
rect 1580 -1253 1660 -1207
rect 1580 -1287 1603 -1253
rect 1637 -1287 1660 -1253
rect 1580 -1333 1660 -1287
rect 1580 -1367 1603 -1333
rect 1637 -1367 1660 -1333
rect 1580 -1413 1660 -1367
rect 1580 -1447 1603 -1413
rect 1637 -1447 1660 -1413
rect 1580 -1480 1660 -1447
rect 1760 -1173 1840 -1080
rect 2300 -1103 2380 -840
rect 2300 -1137 2323 -1103
rect 2357 -1137 2380 -1103
rect 2300 -1170 2380 -1137
rect 2440 -1083 2520 -840
rect 2440 -1117 2463 -1083
rect 2497 -1117 2520 -1083
rect 2440 -1163 2520 -1117
rect 1760 -1207 1783 -1173
rect 1817 -1207 1840 -1173
rect 1760 -1253 1840 -1207
rect 1760 -1287 1783 -1253
rect 1817 -1287 1840 -1253
rect 1760 -1333 1840 -1287
rect 1760 -1367 1783 -1333
rect 1817 -1367 1840 -1333
rect 1760 -1413 1840 -1367
rect 2440 -1197 2463 -1163
rect 2497 -1197 2520 -1163
rect 2440 -1243 2520 -1197
rect 2440 -1277 2463 -1243
rect 2497 -1277 2520 -1243
rect 2440 -1323 2520 -1277
rect 2440 -1357 2463 -1323
rect 2497 -1357 2520 -1323
rect 1760 -1447 1783 -1413
rect 1817 -1447 1840 -1413
rect 750 -1593 950 -1560
rect 750 -1627 783 -1593
rect 817 -1627 883 -1593
rect 917 -1627 950 -1593
rect 750 -1660 950 -1627
rect 1540 -1593 1710 -1560
rect 1540 -1627 1563 -1593
rect 1597 -1627 1653 -1593
rect 1687 -1627 1710 -1593
rect 1540 -1660 1710 -1627
rect -150 -2193 710 -2170
rect -150 -2227 -127 -2193
rect -93 -2227 710 -2193
rect -150 -2250 710 -2227
rect -1510 -2273 -1470 -2270
rect -1510 -2307 -1507 -2273
rect -1473 -2307 -1470 -2273
rect -1510 -2310 -1470 -2307
rect -1430 -2273 -1390 -2270
rect -1430 -2307 -1427 -2273
rect -1393 -2307 -1390 -2273
rect -1430 -2310 -1390 -2307
rect 810 -2330 890 -1660
rect 1760 -2100 1840 -1447
rect 1900 -1423 1980 -1390
rect 1900 -1457 1923 -1423
rect 1957 -1457 1980 -1423
rect 1900 -1490 1980 -1457
rect 2440 -1403 2520 -1357
rect 2440 -1437 2463 -1403
rect 2497 -1437 2520 -1403
rect 2440 -1483 2520 -1437
rect 2440 -1517 2463 -1483
rect 2497 -1517 2520 -1483
rect 2440 -1563 2520 -1517
rect 2440 -1597 2463 -1563
rect 2497 -1597 2520 -1563
rect 2440 -1643 2520 -1597
rect 2440 -1677 2463 -1643
rect 2497 -1677 2520 -1643
rect 2440 -1723 2520 -1677
rect 2440 -1757 2463 -1723
rect 2497 -1757 2520 -1723
rect 2440 -1803 2520 -1757
rect 2440 -1837 2463 -1803
rect 2497 -1837 2520 -1803
rect 2440 -1860 2520 -1837
rect 2620 -1083 2700 -1060
rect 2620 -1117 2643 -1083
rect 2677 -1117 2700 -1083
rect 2620 -1163 2700 -1117
rect 2620 -1197 2643 -1163
rect 2677 -1197 2700 -1163
rect 2620 -1243 2700 -1197
rect 2620 -1277 2643 -1243
rect 2677 -1277 2700 -1243
rect 2620 -1323 2700 -1277
rect 2620 -1357 2643 -1323
rect 2677 -1357 2700 -1323
rect 2620 -1403 2700 -1357
rect 2620 -1437 2643 -1403
rect 2677 -1437 2700 -1403
rect 2620 -1483 2700 -1437
rect 2620 -1517 2643 -1483
rect 2677 -1517 2700 -1483
rect 2620 -1563 2700 -1517
rect 2620 -1597 2643 -1563
rect 2677 -1597 2700 -1563
rect 2620 -1643 2700 -1597
rect 2620 -1677 2643 -1643
rect 2677 -1677 2700 -1643
rect 2620 -1723 2700 -1677
rect 2620 -1757 2643 -1723
rect 2677 -1757 2700 -1723
rect 2620 -1803 2700 -1757
rect 2620 -1837 2643 -1803
rect 2677 -1837 2700 -1803
rect 2520 -1973 2580 -1940
rect 2520 -2007 2533 -1973
rect 2567 -2007 2580 -1973
rect 2520 -2040 2580 -2007
rect 2620 -2100 2700 -1837
rect 2800 -1083 2880 -1060
rect 2800 -1117 2823 -1083
rect 2857 -1117 2880 -1083
rect 2800 -1163 2880 -1117
rect 2800 -1197 2823 -1163
rect 2857 -1197 2880 -1163
rect 2800 -1243 2880 -1197
rect 2800 -1277 2823 -1243
rect 2857 -1277 2880 -1243
rect 2800 -1323 2880 -1277
rect 2800 -1357 2823 -1323
rect 2857 -1357 2880 -1323
rect 2800 -1403 2880 -1357
rect 2800 -1437 2823 -1403
rect 2857 -1437 2880 -1403
rect 2800 -1483 2880 -1437
rect 2800 -1517 2823 -1483
rect 2857 -1517 2880 -1483
rect 2800 -1563 2880 -1517
rect 2800 -1597 2823 -1563
rect 2857 -1597 2880 -1563
rect 2800 -1643 2880 -1597
rect 2800 -1677 2823 -1643
rect 2857 -1677 2880 -1643
rect 2800 -1723 2880 -1677
rect 2800 -1757 2823 -1723
rect 2857 -1757 2880 -1723
rect 2800 -1803 2880 -1757
rect 2800 -1837 2823 -1803
rect 2857 -1837 2880 -1803
rect 2800 -1860 2880 -1837
rect 2740 -1973 2800 -1940
rect 2740 -2007 2753 -1973
rect 2787 -2007 2800 -1973
rect 2740 -2040 2800 -2007
rect 3120 -2100 3220 -10
rect 1760 -2200 3220 -2100
rect -1110 -2363 2880 -2330
rect -1110 -2397 2823 -2363
rect 2857 -2397 2880 -2363
rect -1110 -2430 2880 -2397
rect -1110 -2550 -1010 -2430
rect -1540 -2583 -1010 -2550
rect -1540 -2617 -1507 -2583
rect -1473 -2617 -1010 -2583
rect -1540 -2650 -1010 -2617
rect -400 -2603 570 -2580
rect -400 -2637 -377 -2603
rect -343 -2637 513 -2603
rect 547 -2637 570 -2603
rect -400 -2660 570 -2637
rect -40 -3083 40 -3060
rect -40 -3117 -17 -3083
rect 17 -3117 40 -3083
rect -40 -3140 40 -3117
rect 2630 -3120 2690 -2920
<< viali >>
rect -517 293 -483 327
rect -267 473 -233 507
rect 503 473 537 507
rect 603 473 637 507
rect 233 303 267 337
rect 373 303 407 337
rect -197 143 -163 177
rect -197 63 -163 97
rect 373 223 407 257
rect 553 63 587 97
rect 1563 473 1597 507
rect 1743 473 1777 507
rect 1923 473 1957 507
rect 2663 463 2697 497
rect 733 303 767 337
rect 733 223 767 257
rect 913 63 947 97
rect 1333 303 1367 337
rect 1473 303 1507 337
rect 1473 223 1507 257
rect 1653 63 1687 97
rect 1833 303 1867 337
rect 1833 223 1867 257
rect 2433 293 2467 327
rect 2013 63 2047 97
rect 2573 133 2607 167
rect 2573 53 2607 87
rect -447 -1107 -413 -1073
rect -307 -1107 -273 -1073
rect -307 -1187 -273 -1153
rect -1597 -1557 -1563 -1523
rect -1727 -1977 -1693 -1943
rect -307 -1747 -273 -1713
rect -307 -1827 -273 -1793
rect -1447 -1957 -1413 -1923
rect -237 -1997 -203 -1963
rect 53 -1107 87 -1073
rect 53 -1187 87 -1153
rect 513 -1137 547 -1103
rect 653 -1147 687 -1113
rect 53 -1747 87 -1713
rect 53 -1827 87 -1793
rect 653 -1227 687 -1193
rect -17 -1997 17 -1963
rect 1013 -1147 1047 -1113
rect 1013 -1227 1047 -1193
rect 1423 -1207 1457 -1173
rect 1423 -1287 1457 -1253
rect 2323 -1137 2357 -1103
rect 2463 -1117 2497 -1083
rect 1783 -1207 1817 -1173
rect 1783 -1287 1817 -1253
rect 2463 -1197 2497 -1163
rect 783 -1627 817 -1593
rect 883 -1627 917 -1593
rect 1563 -1627 1597 -1593
rect 1653 -1627 1687 -1593
rect -127 -2227 -93 -2193
rect -1507 -2307 -1473 -2273
rect -1427 -2307 -1393 -2273
rect 1923 -1457 1957 -1423
rect 2463 -1757 2497 -1723
rect 2463 -1837 2497 -1803
rect 2533 -2007 2567 -1973
rect 2823 -1117 2857 -1083
rect 2823 -1197 2857 -1163
rect 2823 -1757 2857 -1723
rect 2823 -1837 2857 -1803
rect 2753 -2007 2787 -1973
rect 2823 -2397 2857 -2363
rect -1507 -2617 -1473 -2583
rect -377 -2637 -343 -2603
rect 513 -2637 547 -2603
rect -17 -3117 17 -3083
<< metal1 >>
rect -320 507 -220 540
rect -320 473 -267 507
rect -233 473 -220 507
rect -320 440 -220 473
rect 430 507 890 540
rect 430 473 503 507
rect 537 473 603 507
rect 637 473 890 507
rect 430 440 890 473
rect 1530 507 1990 540
rect 1530 473 1563 507
rect 1597 473 1743 507
rect 1777 473 1923 507
rect 1957 473 1990 507
rect 1530 440 1990 473
rect 2630 497 2730 530
rect 2630 463 2663 497
rect 2697 463 2730 497
rect 2630 430 2730 463
rect -540 327 -460 360
rect -540 293 -517 327
rect -483 293 -460 327
rect -540 260 -460 293
rect 210 337 290 370
rect 210 303 233 337
rect 267 303 290 337
rect 210 270 290 303
rect 350 337 430 360
rect 350 303 373 337
rect 407 330 430 337
rect 710 337 790 360
rect 710 330 733 337
rect 407 303 733 330
rect 767 303 790 337
rect 350 257 790 303
rect 1310 337 1390 370
rect 1310 303 1333 337
rect 1367 303 1390 337
rect 1310 270 1390 303
rect 1450 340 1530 360
rect 1810 340 1890 360
rect 1450 337 1890 340
rect 1450 303 1473 337
rect 1507 303 1833 337
rect 1867 303 1890 337
rect 350 223 373 257
rect 407 230 733 257
rect 407 223 430 230
rect 350 200 430 223
rect 710 223 733 230
rect 767 223 790 257
rect 710 200 790 223
rect 1450 257 1890 303
rect 1450 223 1473 257
rect 1507 230 1833 257
rect 1507 223 1530 230
rect 1450 200 1530 223
rect 1810 223 1833 230
rect 1867 223 1890 257
rect 1810 200 1890 223
rect 2410 327 2490 360
rect 2410 293 2433 327
rect 2467 293 2490 327
rect -220 177 -140 200
rect -220 143 -197 177
rect -163 143 -140 177
rect -220 97 -140 143
rect -220 63 -197 97
rect -163 63 -140 97
rect -220 -380 -140 63
rect 530 97 970 120
rect 530 63 553 97
rect 587 63 913 97
rect 947 63 970 97
rect 530 20 970 63
rect 530 0 610 20
rect 890 0 970 20
rect 1630 97 2070 120
rect 1630 63 1653 97
rect 1687 63 2013 97
rect 2047 63 2070 97
rect 1630 0 2070 63
rect 2410 -380 2490 293
rect 2550 167 2630 190
rect 2550 133 2573 167
rect 2607 133 2630 167
rect 2550 87 2630 133
rect 2550 53 2573 87
rect 2607 53 2630 87
rect 2550 -380 2630 53
rect -220 -460 2630 -380
rect 230 -930 1310 -830
rect -470 -1073 -390 -1040
rect -470 -1107 -447 -1073
rect -413 -1107 -390 -1073
rect -470 -1140 -390 -1107
rect -330 -1073 -250 -1050
rect -330 -1107 -307 -1073
rect -273 -1080 -250 -1073
rect 30 -1073 110 -1050
rect 30 -1080 53 -1073
rect -273 -1107 53 -1080
rect 87 -1107 110 -1073
rect -330 -1153 110 -1107
rect -330 -1187 -307 -1153
rect -273 -1180 53 -1153
rect -273 -1187 -250 -1180
rect -330 -1210 -250 -1187
rect 30 -1187 53 -1180
rect 87 -1187 110 -1153
rect 30 -1210 110 -1187
rect -1620 -1523 -1540 -1340
rect -1320 -1490 -1220 -1340
rect -1620 -1557 -1597 -1523
rect -1563 -1557 -1540 -1523
rect -1620 -1580 -1540 -1557
rect -330 -1713 -250 -1690
rect -330 -1747 -307 -1713
rect -273 -1720 -250 -1713
rect 30 -1713 110 -1690
rect 30 -1720 53 -1713
rect -273 -1747 53 -1720
rect 87 -1747 110 -1713
rect -330 -1793 110 -1747
rect -330 -1827 -307 -1793
rect -273 -1820 53 -1793
rect -273 -1827 -250 -1820
rect -330 -1850 -250 -1827
rect 30 -1827 53 -1820
rect 87 -1827 110 -1793
rect 30 -1850 110 -1827
rect -1860 -1920 -1760 -1850
rect -1320 -1900 -1220 -1850
rect -1860 -1943 -1660 -1920
rect -1860 -1977 -1727 -1943
rect -1693 -1977 -1660 -1943
rect -1860 -2000 -1660 -1977
rect -1480 -1923 -1220 -1900
rect -1480 -1957 -1447 -1923
rect -1413 -1957 -1220 -1923
rect 230 -1930 330 -930
rect -1480 -1980 -1220 -1957
rect -1860 -2150 -1760 -2000
rect -1320 -2150 -1220 -1980
rect -250 -1963 330 -1930
rect -250 -1997 -237 -1963
rect -203 -1997 -17 -1963
rect 17 -1997 330 -1963
rect -250 -2030 330 -1997
rect 490 -1103 570 -1070
rect 490 -1137 513 -1103
rect 547 -1137 570 -1103
rect 490 -1870 570 -1137
rect 630 -1113 710 -1080
rect 630 -1147 653 -1113
rect 687 -1120 710 -1113
rect 990 -1113 1070 -1080
rect 990 -1120 1013 -1113
rect 687 -1147 1013 -1120
rect 1047 -1147 1070 -1113
rect 630 -1193 1070 -1147
rect 630 -1227 653 -1193
rect 687 -1220 1013 -1193
rect 687 -1227 710 -1220
rect 630 -1250 710 -1227
rect 990 -1227 1013 -1220
rect 1047 -1227 1070 -1193
rect 990 -1250 1070 -1227
rect 1210 -1560 1310 -930
rect 1400 -1173 1480 -1080
rect 1400 -1207 1423 -1173
rect 1457 -1180 1480 -1173
rect 1760 -1173 1840 -1080
rect 2300 -1103 2380 -1070
rect 2300 -1137 2323 -1103
rect 2357 -1137 2380 -1103
rect 2300 -1170 2380 -1137
rect 2440 -1083 2520 -1060
rect 2440 -1117 2463 -1083
rect 2497 -1090 2520 -1083
rect 2800 -1083 2880 -1060
rect 2800 -1090 2823 -1083
rect 2497 -1117 2823 -1090
rect 2857 -1117 2880 -1083
rect 2440 -1163 2880 -1117
rect 1760 -1180 1783 -1173
rect 1457 -1207 1783 -1180
rect 1817 -1207 1840 -1173
rect 1400 -1253 1840 -1207
rect 2440 -1197 2463 -1163
rect 2497 -1190 2823 -1163
rect 2497 -1197 2520 -1190
rect 2440 -1220 2520 -1197
rect 2800 -1197 2823 -1190
rect 2857 -1197 2880 -1163
rect 2800 -1220 2880 -1197
rect 1400 -1287 1423 -1253
rect 1457 -1280 1783 -1253
rect 1457 -1287 1480 -1280
rect 1400 -1310 1480 -1287
rect 1760 -1287 1783 -1280
rect 1817 -1287 1840 -1253
rect 1760 -1310 1840 -1287
rect 1900 -1423 1980 -1390
rect 1900 -1457 1923 -1423
rect 1957 -1457 1980 -1423
rect 710 -1593 990 -1560
rect 710 -1627 783 -1593
rect 817 -1627 883 -1593
rect 917 -1627 990 -1593
rect 710 -1660 990 -1627
rect 1210 -1593 1760 -1560
rect 1210 -1627 1563 -1593
rect 1597 -1627 1653 -1593
rect 1687 -1627 1760 -1593
rect 1210 -1660 1760 -1627
rect 1900 -1870 1980 -1457
rect 2440 -1723 2520 -1700
rect 2440 -1757 2463 -1723
rect 2497 -1730 2520 -1723
rect 2800 -1723 2880 -1700
rect 2800 -1730 2823 -1723
rect 2497 -1757 2823 -1730
rect 2857 -1757 2880 -1723
rect 2440 -1803 2880 -1757
rect 2440 -1837 2463 -1803
rect 2497 -1830 2823 -1803
rect 2497 -1837 2520 -1830
rect 2440 -1860 2520 -1837
rect 2800 -1837 2823 -1830
rect 2857 -1837 2880 -1803
rect 2800 -1860 2880 -1837
rect 490 -1950 1980 -1870
rect -190 -2193 -30 -2140
rect -190 -2227 -127 -2193
rect -93 -2227 -30 -2193
rect -1540 -2273 -1370 -2250
rect -1540 -2307 -1507 -2273
rect -1473 -2307 -1427 -2273
rect -1393 -2307 -1370 -2273
rect -190 -2280 -30 -2227
rect -1540 -2320 -1370 -2307
rect -1850 -3060 -1770 -2390
rect -1540 -2583 -1440 -2320
rect -1540 -2617 -1507 -2583
rect -1473 -2617 -1440 -2583
rect -1540 -2650 -1440 -2617
rect -400 -2603 -320 -2580
rect -400 -2637 -377 -2603
rect -343 -2637 -320 -2603
rect -400 -3060 -320 -2637
rect -150 -2920 -70 -2280
rect 490 -2603 570 -1950
rect 2520 -1973 2880 -1940
rect 2520 -2007 2533 -1973
rect 2567 -2007 2753 -1973
rect 2787 -2007 2880 -1973
rect 2520 -2040 2880 -2007
rect 2800 -2363 2880 -2040
rect 2800 -2397 2823 -2363
rect 2857 -2397 2880 -2363
rect 2800 -2430 2880 -2397
rect 490 -2637 513 -2603
rect 547 -2637 570 -2603
rect 490 -2660 570 -2637
rect -150 -3000 140 -2920
rect -1850 -3083 40 -3060
rect -1850 -3117 -17 -3083
rect 17 -3117 40 -3083
rect -1850 -3140 40 -3117
use sky130_fd_pr__res_xhigh_po_0p35_RSCMUS  sky130_fd_pr__res_xhigh_po_0p35_RSCMUS_0
timestamp 1729593089
transform 0 -1 1378 1 0 -2959
box -191 -1428 191 1428
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0
timestamp 1729593089
transform 0 1 -1812 -1 0 -1488
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1729593089
transform 0 1 -1812 -1 0 -2148
box -38 -48 314 592
<< labels >>
rlabel metal1 s 250 270 250 270 4 B_M3
rlabel locali s 390 0 390 0 4 S1_M3
rlabel locali s 570 0 570 0 4 D1_M3
rlabel locali s 750 0 750 0 4 S2_M3
rlabel locali s 930 0 930 0 4 D2_M3
rlabel poly s 660 -80 660 -80 4 G_M3
rlabel metal1 s 1310 320 1310 320 4 B_M4
rlabel locali s 1490 360 1490 360 4 S1_M4
rlabel locali s 1670 360 1670 360 4 D1_M4
rlabel locali s 1850 360 1850 360 4 S2_M4
rlabel locali s 2030 360 2030 360 4 D2_M4
rlabel metal1 s 1760 540 1760 540 4 G_M4
rlabel metal1 s 2450 360 2450 360 4 B_M2
rlabel locali s 2590 350 2590 350 4 S_M2
rlabel locali s 2770 350 2770 350 4 D_M2
rlabel poly s 2680 -90 2680 -90 4 G_M2
rlabel metal1 s -430 -1140 -430 -1140 4 B_M7
rlabel locali s -290 -1850 -290 -1850 4 S1_M7
rlabel locali s -110 -1850 -110 -1850 4 D_M7
rlabel locali s 70 -1850 70 -1850 4 S2_M7
rlabel metal1 s -110 -2030 -110 -2030 4 G_M7
rlabel metal1 s 2340 -1170 2340 -1170 4 B_M5
rlabel locali s 2660 -1060 2660 -1060 4 D_M5
rlabel locali s 2840 -1860 2840 -1860 4 S2_M5
rlabel metal1 s 2580 -2040 2580 -2040 4 G_M5
rlabel locali s 2480 -1860 2480 -1860 4 S1_M5
rlabel locali s 670 -1080 670 -1080 4 S_M8
rlabel locali s 850 -1480 850 -1480 4 D_M8
rlabel locali s 1030 -1080 1030 -1080 4 S2_M8
rlabel metal1 s 780 -1660 780 -1660 4 G_M8
rlabel metal1 s 1940 -1460 1940 -1460 4 B_M6
rlabel locali s 1800 -1080 1800 -1080 4 S1_M6
rlabel locali s 1620 -1480 1620 -1480 4 D_M6
rlabel locali s 1440 -1080 1440 -1080 4 S2_M6
rlabel metal1 s 1630 -1660 1630 -1660 4 G_M6
rlabel poly s -270 -80 -270 -80 4 G_M1
rlabel locali s -180 360 -180 360 4 D_M1
rlabel locali s -360 0 -360 0 4 S_M1
rlabel metal1 s -500 260 -500 260 4 B_M1
rlabel locali s 1580 -540 1580 -540 4 add_pwr
rlabel metal1 s -110 -2190 -110 -2190 4 input_R
rlabel locali s -1370 -2550 -1370 -2550 4 lock
rlabel locali s -370 740 -370 740 4 VCCA
rlabel metal1 s -1580 -1340 -1580 -1340 4 Dctrl
rlabel metal1 s -270 540 -270 540 4 Vbs1
rlabel metal1 s 2680 530 2680 530 4 Vbs2
rlabel metal1 s 570 540 570 540 4 Vbs3
rlabel metal1 s 1690 540 1690 540 4 Vbs4
rlabel locali s 2930 90 2930 90 4 Isup
rlabel metal1 s -150 -3060 -150 -3060 4 GND
rlabel metal1 s -1270 -1340 -1270 -1340 4 VCCD
<< end >>
