magic
tech sky130A
magscale 1 2
timestamp 1726393621
<< nwell >>
rect -580 -80 -100 440
rect 170 -80 1010 440
rect 1270 -80 2110 440
rect 2370 -90 2850 430
rect -580 -1630 80 -670
rect 2190 -1640 2850 -680
rect 300 -2560 450 -2240
rect 1260 -2250 1430 -2240
rect 1260 -2310 1440 -2250
rect 1260 -2560 1430 -2310
<< pwell >>
rect 380 -1430 1040 -870
rect 1230 -1430 1890 -870
rect 300 -2810 490 -2660
rect 1260 -2810 1470 -2620
<< nmos >>
rect 640 -1350 740 -950
rect 820 -1350 920 -950
rect 1490 -1350 1590 -950
rect 1670 -1350 1770 -950
<< pmoshvt >>
rect -320 0 -220 360
rect 430 0 530 360
rect 610 0 710 360
rect 790 0 890 360
rect 1530 0 1630 360
rect 1710 0 1810 360
rect 1890 0 1990 360
rect 2630 -10 2730 350
rect -320 -1550 -220 -750
rect -140 -1550 -40 -750
rect 2450 -1560 2550 -760
rect 2630 -1560 2730 -760
<< ndiff >>
rect 560 -980 640 -950
rect 560 -1020 580 -980
rect 620 -1020 640 -980
rect 560 -1060 640 -1020
rect 560 -1100 580 -1060
rect 620 -1100 640 -1060
rect 560 -1140 640 -1100
rect 560 -1180 580 -1140
rect 620 -1180 640 -1140
rect 560 -1220 640 -1180
rect 560 -1260 580 -1220
rect 620 -1260 640 -1220
rect 560 -1350 640 -1260
rect 740 -980 820 -950
rect 740 -1020 760 -980
rect 800 -1020 820 -980
rect 740 -1060 820 -1020
rect 740 -1100 760 -1060
rect 800 -1100 820 -1060
rect 740 -1140 820 -1100
rect 740 -1180 760 -1140
rect 800 -1180 820 -1140
rect 740 -1220 820 -1180
rect 740 -1260 760 -1220
rect 800 -1260 820 -1220
rect 740 -1350 820 -1260
rect 920 -980 1000 -950
rect 920 -1020 940 -980
rect 980 -1020 1000 -980
rect 920 -1060 1000 -1020
rect 1410 -980 1490 -950
rect 1410 -1020 1430 -980
rect 1470 -1020 1490 -980
rect 920 -1100 940 -1060
rect 980 -1100 1000 -1060
rect 920 -1140 1000 -1100
rect 920 -1180 940 -1140
rect 980 -1180 1000 -1140
rect 920 -1220 1000 -1180
rect 920 -1260 940 -1220
rect 980 -1260 1000 -1220
rect 920 -1350 1000 -1260
rect 1410 -1060 1490 -1020
rect 1410 -1100 1430 -1060
rect 1470 -1100 1490 -1060
rect 1410 -1140 1490 -1100
rect 1410 -1180 1430 -1140
rect 1470 -1180 1490 -1140
rect 1410 -1220 1490 -1180
rect 1410 -1260 1430 -1220
rect 1470 -1260 1490 -1220
rect 1410 -1350 1490 -1260
rect 1590 -980 1670 -950
rect 1590 -1020 1610 -980
rect 1650 -1020 1670 -980
rect 1590 -1060 1670 -1020
rect 1590 -1100 1610 -1060
rect 1650 -1100 1670 -1060
rect 1590 -1140 1670 -1100
rect 1590 -1180 1610 -1140
rect 1650 -1180 1670 -1140
rect 1590 -1220 1670 -1180
rect 1590 -1260 1610 -1220
rect 1650 -1260 1670 -1220
rect 1590 -1350 1670 -1260
rect 1770 -980 1850 -950
rect 1770 -1020 1790 -980
rect 1830 -1020 1850 -980
rect 1770 -1060 1850 -1020
rect 1770 -1100 1790 -1060
rect 1830 -1100 1850 -1060
rect 1770 -1140 1850 -1100
rect 1770 -1180 1790 -1140
rect 1830 -1180 1850 -1140
rect 1770 -1220 1850 -1180
rect 1770 -1260 1790 -1220
rect 1830 -1260 1850 -1220
rect 1770 -1350 1850 -1260
<< pdiff >>
rect -400 340 -320 360
rect -400 300 -380 340
rect -340 300 -320 340
rect -400 260 -320 300
rect -400 220 -380 260
rect -340 220 -320 260
rect -400 180 -320 220
rect -400 140 -380 180
rect -340 140 -320 180
rect -400 100 -320 140
rect -400 60 -380 100
rect -340 60 -320 100
rect -400 0 -320 60
rect -220 340 -140 360
rect -220 300 -200 340
rect -160 300 -140 340
rect -220 260 -140 300
rect 350 340 430 360
rect 350 300 370 340
rect 410 300 430 340
rect -220 220 -200 260
rect -160 220 -140 260
rect -220 180 -140 220
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 0 -140 60
rect 350 260 430 300
rect 350 220 370 260
rect 410 220 430 260
rect 350 180 430 220
rect 350 140 370 180
rect 410 140 430 180
rect 350 100 430 140
rect 350 60 370 100
rect 410 60 430 100
rect 350 0 430 60
rect 530 340 610 360
rect 530 300 550 340
rect 590 300 610 340
rect 530 260 610 300
rect 530 220 550 260
rect 590 220 610 260
rect 530 180 610 220
rect 530 140 550 180
rect 590 140 610 180
rect 530 100 610 140
rect 530 60 550 100
rect 590 60 610 100
rect 530 0 610 60
rect 710 340 790 360
rect 710 300 730 340
rect 770 300 790 340
rect 710 260 790 300
rect 710 220 730 260
rect 770 220 790 260
rect 710 180 790 220
rect 710 140 730 180
rect 770 140 790 180
rect 710 100 790 140
rect 710 60 730 100
rect 770 60 790 100
rect 710 0 790 60
rect 890 340 970 360
rect 890 300 910 340
rect 950 300 970 340
rect 890 260 970 300
rect 1450 340 1530 360
rect 1450 300 1470 340
rect 1510 300 1530 340
rect 890 220 910 260
rect 950 220 970 260
rect 890 180 970 220
rect 890 140 910 180
rect 950 140 970 180
rect 890 100 970 140
rect 890 60 910 100
rect 950 60 970 100
rect 890 0 970 60
rect 1450 260 1530 300
rect 1450 220 1470 260
rect 1510 220 1530 260
rect 1450 180 1530 220
rect 1450 140 1470 180
rect 1510 140 1530 180
rect 1450 100 1530 140
rect 1450 60 1470 100
rect 1510 60 1530 100
rect 1450 0 1530 60
rect 1630 340 1710 360
rect 1630 300 1650 340
rect 1690 300 1710 340
rect 1630 260 1710 300
rect 1630 220 1650 260
rect 1690 220 1710 260
rect 1630 180 1710 220
rect 1630 140 1650 180
rect 1690 140 1710 180
rect 1630 100 1710 140
rect 1630 60 1650 100
rect 1690 60 1710 100
rect 1630 0 1710 60
rect 1810 340 1890 360
rect 1810 300 1830 340
rect 1870 300 1890 340
rect 1810 260 1890 300
rect 1810 220 1830 260
rect 1870 220 1890 260
rect 1810 180 1890 220
rect 1810 140 1830 180
rect 1870 140 1890 180
rect 1810 100 1890 140
rect 1810 60 1830 100
rect 1870 60 1890 100
rect 1810 0 1890 60
rect 1990 340 2070 360
rect 1990 300 2010 340
rect 2050 300 2070 340
rect 1990 260 2070 300
rect 2550 330 2630 350
rect 2550 290 2570 330
rect 2610 290 2630 330
rect 1990 220 2010 260
rect 2050 220 2070 260
rect 1990 180 2070 220
rect 1990 140 2010 180
rect 2050 140 2070 180
rect 1990 100 2070 140
rect 1990 60 2010 100
rect 2050 60 2070 100
rect 1990 0 2070 60
rect 2550 250 2630 290
rect 2550 210 2570 250
rect 2610 210 2630 250
rect 2550 170 2630 210
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -10 2630 50
rect 2730 330 2810 350
rect 2730 290 2750 330
rect 2790 290 2810 330
rect 2730 250 2810 290
rect 2730 210 2750 250
rect 2790 210 2810 250
rect 2730 170 2810 210
rect 2730 130 2750 170
rect 2790 130 2810 170
rect 2730 90 2810 130
rect 2730 50 2750 90
rect 2790 50 2810 90
rect 2730 -10 2810 50
rect -400 -770 -320 -750
rect -400 -810 -380 -770
rect -340 -810 -320 -770
rect -400 -850 -320 -810
rect -400 -890 -380 -850
rect -340 -890 -320 -850
rect -400 -930 -320 -890
rect -400 -970 -380 -930
rect -340 -970 -320 -930
rect -400 -1010 -320 -970
rect -400 -1050 -380 -1010
rect -340 -1050 -320 -1010
rect -400 -1090 -320 -1050
rect -400 -1130 -380 -1090
rect -340 -1130 -320 -1090
rect -400 -1170 -320 -1130
rect -400 -1210 -380 -1170
rect -340 -1210 -320 -1170
rect -400 -1250 -320 -1210
rect -400 -1290 -380 -1250
rect -340 -1290 -320 -1250
rect -400 -1330 -320 -1290
rect -400 -1370 -380 -1330
rect -340 -1370 -320 -1330
rect -400 -1410 -320 -1370
rect -400 -1450 -380 -1410
rect -340 -1450 -320 -1410
rect -400 -1490 -320 -1450
rect -400 -1530 -380 -1490
rect -340 -1530 -320 -1490
rect -400 -1550 -320 -1530
rect -220 -770 -140 -750
rect -220 -810 -200 -770
rect -160 -810 -140 -770
rect -220 -850 -140 -810
rect -220 -890 -200 -850
rect -160 -890 -140 -850
rect -220 -930 -140 -890
rect -220 -970 -200 -930
rect -160 -970 -140 -930
rect -220 -1010 -140 -970
rect -220 -1050 -200 -1010
rect -160 -1050 -140 -1010
rect -220 -1090 -140 -1050
rect -220 -1130 -200 -1090
rect -160 -1130 -140 -1090
rect -220 -1170 -140 -1130
rect -220 -1210 -200 -1170
rect -160 -1210 -140 -1170
rect -220 -1250 -140 -1210
rect -220 -1290 -200 -1250
rect -160 -1290 -140 -1250
rect -220 -1330 -140 -1290
rect -220 -1370 -200 -1330
rect -160 -1370 -140 -1330
rect -220 -1410 -140 -1370
rect -220 -1450 -200 -1410
rect -160 -1450 -140 -1410
rect -220 -1490 -140 -1450
rect -220 -1530 -200 -1490
rect -160 -1530 -140 -1490
rect -220 -1550 -140 -1530
rect -40 -770 40 -750
rect -40 -810 -20 -770
rect 20 -810 40 -770
rect -40 -850 40 -810
rect -40 -890 -20 -850
rect 20 -890 40 -850
rect 2370 -780 2450 -760
rect 2370 -820 2390 -780
rect 2430 -820 2450 -780
rect 2370 -860 2450 -820
rect -40 -930 40 -890
rect -40 -970 -20 -930
rect 20 -970 40 -930
rect -40 -1010 40 -970
rect -40 -1050 -20 -1010
rect 20 -1050 40 -1010
rect -40 -1090 40 -1050
rect -40 -1130 -20 -1090
rect 20 -1130 40 -1090
rect -40 -1170 40 -1130
rect -40 -1210 -20 -1170
rect 20 -1210 40 -1170
rect -40 -1250 40 -1210
rect -40 -1290 -20 -1250
rect 20 -1290 40 -1250
rect -40 -1330 40 -1290
rect -40 -1370 -20 -1330
rect 20 -1370 40 -1330
rect 2370 -900 2390 -860
rect 2430 -900 2450 -860
rect 2370 -940 2450 -900
rect 2370 -980 2390 -940
rect 2430 -980 2450 -940
rect 2370 -1020 2450 -980
rect 2370 -1060 2390 -1020
rect 2430 -1060 2450 -1020
rect 2370 -1100 2450 -1060
rect 2370 -1140 2390 -1100
rect 2430 -1140 2450 -1100
rect 2370 -1180 2450 -1140
rect 2370 -1220 2390 -1180
rect 2430 -1220 2450 -1180
rect 2370 -1260 2450 -1220
rect 2370 -1300 2390 -1260
rect 2430 -1300 2450 -1260
rect 2370 -1340 2450 -1300
rect -40 -1410 40 -1370
rect -40 -1450 -20 -1410
rect 20 -1450 40 -1410
rect -40 -1490 40 -1450
rect -40 -1530 -20 -1490
rect 20 -1530 40 -1490
rect 2370 -1380 2390 -1340
rect 2430 -1380 2450 -1340
rect 2370 -1420 2450 -1380
rect 2370 -1460 2390 -1420
rect 2430 -1460 2450 -1420
rect 2370 -1500 2450 -1460
rect -40 -1550 40 -1530
rect 2370 -1540 2390 -1500
rect 2430 -1540 2450 -1500
rect 2370 -1560 2450 -1540
rect 2550 -780 2630 -760
rect 2550 -820 2570 -780
rect 2610 -820 2630 -780
rect 2550 -860 2630 -820
rect 2550 -900 2570 -860
rect 2610 -900 2630 -860
rect 2550 -940 2630 -900
rect 2550 -980 2570 -940
rect 2610 -980 2630 -940
rect 2550 -1020 2630 -980
rect 2550 -1060 2570 -1020
rect 2610 -1060 2630 -1020
rect 2550 -1100 2630 -1060
rect 2550 -1140 2570 -1100
rect 2610 -1140 2630 -1100
rect 2550 -1180 2630 -1140
rect 2550 -1220 2570 -1180
rect 2610 -1220 2630 -1180
rect 2550 -1260 2630 -1220
rect 2550 -1300 2570 -1260
rect 2610 -1300 2630 -1260
rect 2550 -1340 2630 -1300
rect 2550 -1380 2570 -1340
rect 2610 -1380 2630 -1340
rect 2550 -1420 2630 -1380
rect 2550 -1460 2570 -1420
rect 2610 -1460 2630 -1420
rect 2550 -1500 2630 -1460
rect 2550 -1540 2570 -1500
rect 2610 -1540 2630 -1500
rect 2550 -1560 2630 -1540
rect 2730 -780 2810 -760
rect 2730 -820 2750 -780
rect 2790 -820 2810 -780
rect 2730 -860 2810 -820
rect 2730 -900 2750 -860
rect 2790 -900 2810 -860
rect 2730 -940 2810 -900
rect 2730 -980 2750 -940
rect 2790 -980 2810 -940
rect 2730 -1020 2810 -980
rect 2730 -1060 2750 -1020
rect 2790 -1060 2810 -1020
rect 2730 -1100 2810 -1060
rect 2730 -1140 2750 -1100
rect 2790 -1140 2810 -1100
rect 2730 -1180 2810 -1140
rect 2730 -1220 2750 -1180
rect 2790 -1220 2810 -1180
rect 2730 -1260 2810 -1220
rect 2730 -1300 2750 -1260
rect 2790 -1300 2810 -1260
rect 2730 -1340 2810 -1300
rect 2730 -1380 2750 -1340
rect 2790 -1380 2810 -1340
rect 2730 -1420 2810 -1380
rect 2730 -1460 2750 -1420
rect 2790 -1460 2810 -1420
rect 2730 -1500 2810 -1460
rect 2730 -1540 2750 -1500
rect 2790 -1540 2810 -1500
rect 2730 -1560 2810 -1540
<< ndiffc >>
rect 580 -1020 620 -980
rect 580 -1100 620 -1060
rect 580 -1180 620 -1140
rect 580 -1260 620 -1220
rect 760 -1020 800 -980
rect 760 -1100 800 -1060
rect 760 -1180 800 -1140
rect 760 -1260 800 -1220
rect 940 -1020 980 -980
rect 1430 -1020 1470 -980
rect 940 -1100 980 -1060
rect 940 -1180 980 -1140
rect 940 -1260 980 -1220
rect 1430 -1100 1470 -1060
rect 1430 -1180 1470 -1140
rect 1430 -1260 1470 -1220
rect 1610 -1020 1650 -980
rect 1610 -1100 1650 -1060
rect 1610 -1180 1650 -1140
rect 1610 -1260 1650 -1220
rect 1790 -1020 1830 -980
rect 1790 -1100 1830 -1060
rect 1790 -1180 1830 -1140
rect 1790 -1260 1830 -1220
<< pdiffc >>
rect -380 300 -340 340
rect -380 220 -340 260
rect -380 140 -340 180
rect -380 60 -340 100
rect -200 300 -160 340
rect 370 300 410 340
rect -200 220 -160 260
rect -200 140 -160 180
rect -200 60 -160 100
rect 370 220 410 260
rect 370 140 410 180
rect 370 60 410 100
rect 550 300 590 340
rect 550 220 590 260
rect 550 140 590 180
rect 550 60 590 100
rect 730 300 770 340
rect 730 220 770 260
rect 730 140 770 180
rect 730 60 770 100
rect 910 300 950 340
rect 1470 300 1510 340
rect 910 220 950 260
rect 910 140 950 180
rect 910 60 950 100
rect 1470 220 1510 260
rect 1470 140 1510 180
rect 1470 60 1510 100
rect 1650 300 1690 340
rect 1650 220 1690 260
rect 1650 140 1690 180
rect 1650 60 1690 100
rect 1830 300 1870 340
rect 1830 220 1870 260
rect 1830 140 1870 180
rect 1830 60 1870 100
rect 2010 300 2050 340
rect 2570 290 2610 330
rect 2010 220 2050 260
rect 2010 140 2050 180
rect 2010 60 2050 100
rect 2570 210 2610 250
rect 2570 130 2610 170
rect 2570 50 2610 90
rect 2750 290 2790 330
rect 2750 210 2790 250
rect 2750 130 2790 170
rect 2750 50 2790 90
rect -380 -810 -340 -770
rect -380 -890 -340 -850
rect -380 -970 -340 -930
rect -380 -1050 -340 -1010
rect -380 -1130 -340 -1090
rect -380 -1210 -340 -1170
rect -380 -1290 -340 -1250
rect -380 -1370 -340 -1330
rect -380 -1450 -340 -1410
rect -380 -1530 -340 -1490
rect -200 -810 -160 -770
rect -200 -890 -160 -850
rect -200 -970 -160 -930
rect -200 -1050 -160 -1010
rect -200 -1130 -160 -1090
rect -200 -1210 -160 -1170
rect -200 -1290 -160 -1250
rect -200 -1370 -160 -1330
rect -200 -1450 -160 -1410
rect -200 -1530 -160 -1490
rect -20 -810 20 -770
rect -20 -890 20 -850
rect 2390 -820 2430 -780
rect -20 -970 20 -930
rect -20 -1050 20 -1010
rect -20 -1130 20 -1090
rect -20 -1210 20 -1170
rect -20 -1290 20 -1250
rect -20 -1370 20 -1330
rect 2390 -900 2430 -860
rect 2390 -980 2430 -940
rect 2390 -1060 2430 -1020
rect 2390 -1140 2430 -1100
rect 2390 -1220 2430 -1180
rect 2390 -1300 2430 -1260
rect -20 -1450 20 -1410
rect -20 -1530 20 -1490
rect 2390 -1380 2430 -1340
rect 2390 -1460 2430 -1420
rect 2390 -1540 2430 -1500
rect 2570 -820 2610 -780
rect 2570 -900 2610 -860
rect 2570 -980 2610 -940
rect 2570 -1060 2610 -1020
rect 2570 -1140 2610 -1100
rect 2570 -1220 2610 -1180
rect 2570 -1300 2610 -1260
rect 2570 -1380 2610 -1340
rect 2570 -1460 2610 -1420
rect 2570 -1540 2610 -1500
rect 2750 -820 2790 -780
rect 2750 -900 2790 -860
rect 2750 -980 2790 -940
rect 2750 -1060 2790 -1020
rect 2750 -1140 2790 -1100
rect 2750 -1220 2790 -1180
rect 2750 -1300 2790 -1260
rect 2750 -1380 2790 -1340
rect 2750 -1460 2790 -1420
rect 2750 -1540 2790 -1500
<< psubdiff >>
rect 420 -970 500 -940
rect 420 -1010 440 -970
rect 480 -1010 500 -970
rect 420 -1040 500 -1010
rect 1270 -970 1350 -940
rect 1270 -1010 1290 -970
rect 1330 -1010 1350 -970
rect 1270 -1040 1350 -1010
rect 1300 -2690 1380 -2660
rect 340 -2720 420 -2690
rect 340 -2760 360 -2720
rect 400 -2760 420 -2720
rect 1300 -2730 1320 -2690
rect 1360 -2730 1380 -2690
rect 1300 -2760 1380 -2730
rect 340 -2790 420 -2760
<< nsubdiff >>
rect -540 330 -460 360
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect 210 340 290 370
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 1310 270 1390 300
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect 2410 260 2490 290
rect -540 -770 -460 -740
rect -540 -810 -520 -770
rect -480 -810 -460 -770
rect -540 -840 -460 -810
rect 2230 -800 2310 -770
rect 2230 -840 2250 -800
rect 2290 -840 2310 -800
rect 2230 -870 2310 -840
rect 340 -2380 420 -2350
rect 340 -2420 360 -2380
rect 400 -2420 420 -2380
rect 340 -2450 420 -2420
rect 1300 -2380 1380 -2350
rect 1300 -2420 1320 -2380
rect 1360 -2420 1380 -2380
rect 1300 -2450 1380 -2420
<< psubdiffcont >>
rect 440 -1010 480 -970
rect 1290 -1010 1330 -970
rect 360 -2760 400 -2720
rect 1320 -2730 1360 -2690
<< nsubdiffcont >>
rect -520 290 -480 330
rect 230 300 270 340
rect 1330 300 1370 340
rect 2430 290 2470 330
rect -520 -810 -480 -770
rect 2250 -840 2290 -800
rect 360 -2420 400 -2380
rect 1320 -2420 1360 -2380
<< poly >>
rect -320 510 -220 540
rect -320 470 -270 510
rect -230 470 -220 510
rect -320 360 -220 470
rect 430 510 890 540
rect 430 470 500 510
rect 540 470 600 510
rect 640 470 890 510
rect 430 440 890 470
rect 430 360 530 440
rect 610 360 710 440
rect 790 360 890 440
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 1530 360 1630 440
rect 1710 360 1810 440
rect 1890 360 1990 440
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 350 2730 460
rect -320 -80 -220 0
rect 430 -80 530 0
rect 610 -80 710 0
rect 790 -80 890 0
rect 1530 -80 1630 0
rect 1710 -80 1810 0
rect 1890 -80 1990 0
rect 2630 -90 2730 -10
rect -320 -750 -220 -670
rect -140 -750 -40 -670
rect 2450 -760 2550 -680
rect 2630 -760 2730 -680
rect 1490 -800 1770 -770
rect 1490 -840 1500 -800
rect 1540 -840 1720 -800
rect 1760 -840 1770 -800
rect 1490 -870 1770 -840
rect 640 -950 740 -870
rect 820 -950 920 -870
rect 1490 -950 1590 -870
rect 1670 -950 1770 -870
rect 640 -1430 740 -1350
rect 820 -1430 920 -1350
rect 1490 -1430 1590 -1350
rect 1670 -1430 1770 -1350
rect 640 -1460 920 -1430
rect 640 -1500 710 -1460
rect 750 -1500 810 -1460
rect 850 -1500 920 -1460
rect 640 -1530 920 -1500
rect -320 -1630 -220 -1550
rect -140 -1630 -40 -1550
rect -320 -1660 -40 -1630
rect -320 -1700 -310 -1660
rect -270 -1700 -90 -1660
rect -50 -1700 -40 -1660
rect -320 -1730 -40 -1700
rect 2450 -1640 2550 -1560
rect 2630 -1640 2730 -1560
rect 2450 -1670 2730 -1640
rect 2450 -1710 2460 -1670
rect 2500 -1710 2680 -1670
rect 2720 -1710 2730 -1670
rect 2450 -1740 2730 -1710
<< polycont >>
rect -270 470 -230 510
rect 500 470 540 510
rect 600 470 640 510
rect 1560 470 1600 510
rect 1740 470 1780 510
rect 1920 470 1960 510
rect 2660 460 2700 500
rect 1500 -840 1540 -800
rect 1720 -840 1760 -800
rect 710 -1500 750 -1460
rect 810 -1500 850 -1460
rect -310 -1700 -270 -1660
rect -90 -1700 -50 -1660
rect 2460 -1710 2500 -1670
rect 2680 -1710 2720 -1670
<< locali >>
rect -540 740 790 840
rect -540 330 -460 740
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect -400 340 -320 740
rect -280 510 -220 540
rect -280 470 -270 510
rect -230 470 -220 510
rect -280 440 -220 470
rect -400 300 -380 340
rect -340 300 -320 340
rect -400 260 -320 300
rect -400 220 -380 260
rect -340 220 -320 260
rect -400 180 -320 220
rect -400 140 -380 180
rect -340 140 -320 180
rect -400 100 -320 140
rect -400 60 -380 100
rect -340 60 -320 100
rect -400 0 -320 60
rect -220 340 -140 360
rect -220 300 -200 340
rect -160 300 -140 340
rect -220 260 -140 300
rect 210 340 290 740
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 350 340 430 740
rect 470 510 670 540
rect 470 470 500 510
rect 540 470 600 510
rect 640 470 670 510
rect 470 440 670 470
rect 350 300 370 340
rect 410 300 430 340
rect -220 220 -200 260
rect -160 220 -140 260
rect -220 180 -140 220
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 0 -140 60
rect 350 260 430 300
rect 350 220 370 260
rect 410 220 430 260
rect 350 180 430 220
rect 350 140 370 180
rect 410 140 430 180
rect 350 100 430 140
rect 350 60 370 100
rect 410 60 430 100
rect 350 0 430 60
rect 530 340 610 360
rect 530 300 550 340
rect 590 300 610 340
rect 530 260 610 300
rect 530 220 550 260
rect 590 220 610 260
rect 530 180 610 220
rect 530 140 550 180
rect 590 140 610 180
rect 530 100 610 140
rect 530 60 550 100
rect 590 60 610 100
rect 530 0 610 60
rect 710 340 790 740
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 430 2730 460
rect 710 300 730 340
rect 770 300 790 340
rect 710 260 790 300
rect 710 220 730 260
rect 770 220 790 260
rect 710 180 790 220
rect 710 140 730 180
rect 770 140 790 180
rect 710 100 790 140
rect 710 60 730 100
rect 770 60 790 100
rect 710 0 790 60
rect 890 340 970 360
rect 890 300 910 340
rect 950 300 970 340
rect 890 260 970 300
rect 890 220 910 260
rect 950 220 970 260
rect 890 200 970 220
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 1310 200 1390 300
rect 1450 340 1530 360
rect 1450 300 1470 340
rect 1510 300 1530 340
rect 1450 260 1530 300
rect 1450 220 1470 260
rect 1510 220 1530 260
rect 1450 200 1530 220
rect 890 180 1530 200
rect 890 140 910 180
rect 950 140 1470 180
rect 1510 140 1530 180
rect 890 120 1530 140
rect 890 100 970 120
rect 890 60 910 100
rect 950 60 970 100
rect 890 0 970 60
rect 1450 100 1530 120
rect 1450 60 1470 100
rect 1510 60 1530 100
rect 1450 0 1530 60
rect 1630 340 1710 360
rect 1630 300 1650 340
rect 1690 300 1710 340
rect 1630 260 1710 300
rect 1630 220 1650 260
rect 1690 220 1710 260
rect 1630 180 1710 220
rect 1630 140 1650 180
rect 1690 140 1710 180
rect 1630 100 1710 140
rect 1630 60 1650 100
rect 1690 60 1710 100
rect 1630 -440 1710 60
rect 1810 340 1890 360
rect 1810 300 1830 340
rect 1870 300 1890 340
rect 1810 260 1890 300
rect 1810 220 1830 260
rect 1870 220 1890 260
rect 1810 180 1890 220
rect 1810 140 1830 180
rect 1870 140 1890 180
rect 1810 100 1890 140
rect 1810 60 1830 100
rect 1870 60 1890 100
rect 1810 0 1890 60
rect 1990 340 2070 360
rect 1990 300 2010 340
rect 2050 300 2070 340
rect 1990 260 2070 300
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect 2410 260 2490 290
rect 2550 330 2630 350
rect 2550 290 2570 330
rect 2610 290 2630 330
rect 1990 220 2010 260
rect 2050 220 2070 260
rect 1990 180 2070 220
rect 1990 140 2010 180
rect 2050 140 2070 180
rect 1990 100 2070 140
rect 1990 60 2010 100
rect 2050 60 2070 100
rect 1990 -440 2070 60
rect 2550 250 2630 290
rect 2550 210 2570 250
rect 2610 210 2630 250
rect 2550 170 2630 210
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -10 2630 50
rect 2730 330 2810 350
rect 2730 290 2750 330
rect 2790 290 2810 330
rect 2730 250 2810 290
rect 2730 210 2750 250
rect 2790 210 2810 250
rect 2730 170 2810 210
rect 2730 130 2750 170
rect 2790 130 2810 170
rect 2730 90 2810 130
rect 2730 50 2750 90
rect 2790 50 3050 90
rect 2730 -10 3050 50
rect -540 -540 2810 -440
rect -540 -770 -460 -540
rect -540 -810 -520 -770
rect -480 -810 -460 -770
rect -540 -840 -460 -810
rect -400 -770 -320 -540
rect -400 -810 -380 -770
rect -340 -810 -320 -770
rect -400 -850 -320 -810
rect -400 -890 -380 -850
rect -340 -890 -320 -850
rect -400 -930 -320 -890
rect -400 -970 -380 -930
rect -340 -970 -320 -930
rect -400 -1010 -320 -970
rect -400 -1050 -380 -1010
rect -340 -1050 -320 -1010
rect -400 -1090 -320 -1050
rect -400 -1130 -380 -1090
rect -340 -1130 -320 -1090
rect -400 -1170 -320 -1130
rect -400 -1210 -380 -1170
rect -340 -1210 -320 -1170
rect -400 -1250 -320 -1210
rect -400 -1290 -380 -1250
rect -340 -1290 -320 -1250
rect -400 -1330 -320 -1290
rect -400 -1370 -380 -1330
rect -340 -1370 -320 -1330
rect -400 -1410 -320 -1370
rect -400 -1450 -380 -1410
rect -340 -1450 -320 -1410
rect -400 -1490 -320 -1450
rect -400 -1530 -380 -1490
rect -340 -1530 -320 -1490
rect -400 -1550 -320 -1530
rect -220 -770 -140 -750
rect -220 -810 -200 -770
rect -160 -810 -140 -770
rect -220 -850 -140 -810
rect -220 -890 -200 -850
rect -160 -890 -140 -850
rect -220 -930 -140 -890
rect -220 -970 -200 -930
rect -160 -970 -140 -930
rect -220 -1010 -140 -970
rect -220 -1050 -200 -1010
rect -160 -1050 -140 -1010
rect -220 -1090 -140 -1050
rect -220 -1130 -200 -1090
rect -160 -1130 -140 -1090
rect -220 -1170 -140 -1130
rect -220 -1210 -200 -1170
rect -160 -1210 -140 -1170
rect -220 -1250 -140 -1210
rect -220 -1290 -200 -1250
rect -160 -1290 -140 -1250
rect -220 -1330 -140 -1290
rect -220 -1370 -200 -1330
rect -160 -1370 -140 -1330
rect -220 -1410 -140 -1370
rect -220 -1450 -200 -1410
rect -160 -1450 -140 -1410
rect -220 -1490 -140 -1450
rect -220 -1530 -200 -1490
rect -160 -1530 -140 -1490
rect -320 -1660 -260 -1630
rect -320 -1700 -310 -1660
rect -270 -1700 -260 -1660
rect -320 -1730 -260 -1700
rect -220 -1830 -140 -1530
rect -40 -770 40 -540
rect -40 -810 -20 -770
rect 20 -810 40 -770
rect -40 -850 40 -810
rect -40 -890 -20 -850
rect 20 -890 40 -850
rect -40 -930 40 -890
rect -40 -970 -20 -930
rect 20 -970 40 -930
rect -40 -1010 40 -970
rect -40 -1050 -20 -1010
rect 20 -1050 40 -1010
rect -40 -1090 40 -1050
rect -40 -1130 -20 -1090
rect 20 -1130 40 -1090
rect -40 -1170 40 -1130
rect -40 -1210 -20 -1170
rect 20 -1210 40 -1170
rect -40 -1250 40 -1210
rect -40 -1290 -20 -1250
rect 20 -1290 40 -1250
rect -40 -1330 40 -1290
rect -40 -1370 -20 -1330
rect 20 -1370 40 -1330
rect -40 -1410 40 -1370
rect -40 -1450 -20 -1410
rect 20 -1450 40 -1410
rect -40 -1490 40 -1450
rect -40 -1530 -20 -1490
rect 20 -1530 40 -1490
rect -40 -1550 40 -1530
rect 420 -970 500 -940
rect 420 -1010 440 -970
rect 480 -1010 500 -970
rect -100 -1660 -40 -1630
rect -100 -1700 -90 -1660
rect -50 -1700 -40 -1660
rect -100 -1730 -40 -1700
rect 420 -1830 500 -1010
rect 560 -980 640 -950
rect 560 -1020 580 -980
rect 620 -1020 640 -980
rect 560 -1060 640 -1020
rect 560 -1100 580 -1060
rect 620 -1100 640 -1060
rect 560 -1140 640 -1100
rect 560 -1180 580 -1140
rect 620 -1180 640 -1140
rect 560 -1220 640 -1180
rect 560 -1260 580 -1220
rect 620 -1260 640 -1220
rect 560 -1830 640 -1260
rect 740 -980 820 -540
rect 1490 -800 1550 -770
rect 1490 -840 1500 -800
rect 1540 -840 1550 -800
rect 1490 -870 1550 -840
rect 740 -1020 760 -980
rect 800 -1020 820 -980
rect 740 -1060 820 -1020
rect 740 -1100 760 -1060
rect 800 -1100 820 -1060
rect 740 -1140 820 -1100
rect 740 -1180 760 -1140
rect 800 -1180 820 -1140
rect 740 -1220 820 -1180
rect 740 -1260 760 -1220
rect 800 -1260 820 -1220
rect 740 -1350 820 -1260
rect 920 -980 1000 -950
rect 920 -1020 940 -980
rect 980 -1020 1000 -980
rect 920 -1060 1000 -1020
rect 920 -1100 940 -1060
rect 980 -1100 1000 -1060
rect 920 -1140 1000 -1100
rect 920 -1180 940 -1140
rect 980 -1180 1000 -1140
rect 920 -1220 1000 -1180
rect 920 -1260 940 -1220
rect 980 -1260 1000 -1220
rect 680 -1460 880 -1430
rect 680 -1500 710 -1460
rect 750 -1500 810 -1460
rect 850 -1500 880 -1460
rect 680 -1530 880 -1500
rect 920 -1830 1000 -1260
rect -220 -1930 1000 -1830
rect 1270 -970 1350 -940
rect 1270 -1010 1290 -970
rect 1330 -1010 1350 -970
rect 1270 -1830 1350 -1010
rect 1410 -980 1490 -950
rect 1410 -1020 1430 -980
rect 1470 -1020 1490 -980
rect 1410 -1060 1490 -1020
rect 1410 -1100 1430 -1060
rect 1470 -1100 1490 -1060
rect 1410 -1140 1490 -1100
rect 1410 -1180 1430 -1140
rect 1470 -1180 1490 -1140
rect 1410 -1220 1490 -1180
rect 1410 -1260 1430 -1220
rect 1470 -1260 1490 -1220
rect 1410 -1830 1490 -1260
rect 1590 -980 1670 -540
rect 1710 -800 1770 -770
rect 1710 -840 1720 -800
rect 1760 -840 1770 -800
rect 1710 -870 1770 -840
rect 2230 -800 2310 -540
rect 2230 -840 2250 -800
rect 2290 -840 2310 -800
rect 2230 -870 2310 -840
rect 2370 -780 2450 -540
rect 2370 -820 2390 -780
rect 2430 -820 2450 -780
rect 2370 -860 2450 -820
rect 2370 -900 2390 -860
rect 2430 -900 2450 -860
rect 2370 -940 2450 -900
rect 1590 -1020 1610 -980
rect 1650 -1020 1670 -980
rect 1590 -1060 1670 -1020
rect 1590 -1100 1610 -1060
rect 1650 -1100 1670 -1060
rect 1590 -1140 1670 -1100
rect 1590 -1180 1610 -1140
rect 1650 -1180 1670 -1140
rect 1590 -1220 1670 -1180
rect 1590 -1260 1610 -1220
rect 1650 -1260 1670 -1220
rect 1590 -1350 1670 -1260
rect 1770 -980 1850 -950
rect 1770 -1020 1790 -980
rect 1830 -1020 1850 -980
rect 1770 -1060 1850 -1020
rect 1770 -1100 1790 -1060
rect 1830 -1100 1850 -1060
rect 1770 -1140 1850 -1100
rect 1770 -1180 1790 -1140
rect 1830 -1180 1850 -1140
rect 1770 -1220 1850 -1180
rect 1770 -1260 1790 -1220
rect 1830 -1260 1850 -1220
rect 1770 -1830 1850 -1260
rect 2370 -980 2390 -940
rect 2430 -980 2450 -940
rect 2370 -1020 2450 -980
rect 2370 -1060 2390 -1020
rect 2430 -1060 2450 -1020
rect 2370 -1100 2450 -1060
rect 2370 -1140 2390 -1100
rect 2430 -1140 2450 -1100
rect 2370 -1180 2450 -1140
rect 2370 -1220 2390 -1180
rect 2430 -1220 2450 -1180
rect 2370 -1260 2450 -1220
rect 2370 -1300 2390 -1260
rect 2430 -1300 2450 -1260
rect 2370 -1340 2450 -1300
rect 2370 -1380 2390 -1340
rect 2430 -1380 2450 -1340
rect 2370 -1420 2450 -1380
rect 2370 -1460 2390 -1420
rect 2430 -1460 2450 -1420
rect 2370 -1500 2450 -1460
rect 2370 -1540 2390 -1500
rect 2430 -1540 2450 -1500
rect 2370 -1560 2450 -1540
rect 2550 -780 2630 -760
rect 2550 -820 2570 -780
rect 2610 -820 2630 -780
rect 2550 -860 2630 -820
rect 2550 -900 2570 -860
rect 2610 -900 2630 -860
rect 2550 -940 2630 -900
rect 2550 -980 2570 -940
rect 2610 -980 2630 -940
rect 2550 -1020 2630 -980
rect 2550 -1060 2570 -1020
rect 2610 -1060 2630 -1020
rect 2550 -1100 2630 -1060
rect 2550 -1140 2570 -1100
rect 2610 -1140 2630 -1100
rect 2550 -1180 2630 -1140
rect 2550 -1220 2570 -1180
rect 2610 -1220 2630 -1180
rect 2550 -1260 2630 -1220
rect 2550 -1300 2570 -1260
rect 2610 -1300 2630 -1260
rect 2550 -1340 2630 -1300
rect 2550 -1380 2570 -1340
rect 2610 -1380 2630 -1340
rect 2550 -1420 2630 -1380
rect 2550 -1460 2570 -1420
rect 2610 -1460 2630 -1420
rect 2550 -1500 2630 -1460
rect 2550 -1540 2570 -1500
rect 2610 -1540 2630 -1500
rect 2450 -1670 2510 -1640
rect 2450 -1710 2460 -1670
rect 2500 -1710 2510 -1670
rect 2450 -1740 2510 -1710
rect 2550 -1830 2630 -1540
rect 2730 -780 2810 -540
rect 2730 -820 2750 -780
rect 2790 -820 2810 -780
rect 2730 -860 2810 -820
rect 2730 -900 2750 -860
rect 2790 -900 2810 -860
rect 2730 -940 2810 -900
rect 2730 -980 2750 -940
rect 2790 -980 2810 -940
rect 2730 -1020 2810 -980
rect 2730 -1060 2750 -1020
rect 2790 -1060 2810 -1020
rect 2730 -1100 2810 -1060
rect 2730 -1140 2750 -1100
rect 2790 -1140 2810 -1100
rect 2730 -1180 2810 -1140
rect 2730 -1220 2750 -1180
rect 2790 -1220 2810 -1180
rect 2730 -1260 2810 -1220
rect 2730 -1300 2750 -1260
rect 2790 -1300 2810 -1260
rect 2730 -1340 2810 -1300
rect 2730 -1380 2750 -1340
rect 2790 -1380 2810 -1340
rect 2730 -1420 2810 -1380
rect 2730 -1460 2750 -1420
rect 2790 -1460 2810 -1420
rect 2730 -1500 2810 -1460
rect 2730 -1540 2750 -1500
rect 2790 -1540 2810 -1500
rect 2730 -1560 2810 -1540
rect 2670 -1670 2730 -1640
rect 2670 -1710 2680 -1670
rect 2720 -1710 2730 -1670
rect 2670 -1740 2730 -1710
rect 2950 -1830 3050 -10
rect 1270 -1930 3050 -1830
rect -220 -3200 -140 -1930
rect 340 -2380 420 -2350
rect 340 -2420 360 -2380
rect 400 -2420 420 -2380
rect 340 -2450 420 -2420
rect 1300 -2380 1380 -2350
rect 1300 -2420 1320 -2380
rect 1360 -2420 1380 -2380
rect 1300 -2450 1380 -2420
rect 1300 -2690 1380 -2660
rect 340 -2720 420 -2690
rect 340 -2760 360 -2720
rect 400 -2760 420 -2720
rect 1300 -2730 1320 -2690
rect 1360 -2730 1380 -2690
rect 340 -2790 420 -2760
rect -220 -3240 -200 -3200
rect -160 -3240 -140 -3200
rect -220 -3260 -140 -3240
<< viali >>
rect -520 290 -480 330
rect -270 470 -230 510
rect 230 300 270 340
rect 500 470 540 510
rect 600 470 640 510
rect -200 140 -160 180
rect -200 60 -160 100
rect 550 220 590 260
rect 550 140 590 180
rect 550 60 590 100
rect 1560 470 1600 510
rect 1740 470 1780 510
rect 1920 470 1960 510
rect 2660 460 2700 500
rect 910 220 950 260
rect 1330 300 1370 340
rect 1470 220 1510 260
rect 910 140 950 180
rect 1470 140 1510 180
rect 910 60 950 100
rect 1470 60 1510 100
rect 1830 220 1870 260
rect 1830 140 1870 180
rect 1830 60 1870 100
rect 2430 290 2470 330
rect 2570 130 2610 170
rect 2570 50 2610 90
rect -520 -810 -480 -770
rect -310 -1700 -270 -1660
rect 440 -1010 480 -970
rect -90 -1700 -50 -1660
rect 1500 -840 1540 -800
rect 710 -1500 750 -1460
rect 810 -1500 850 -1460
rect 1290 -1010 1330 -970
rect 1720 -840 1760 -800
rect 2460 -1710 2500 -1670
rect 2680 -1710 2720 -1670
rect 360 -2420 400 -2380
rect 1320 -2420 1360 -2380
rect 696 -2478 736 -2438
rect 1580 -2480 1620 -2440
rect 520 -2600 560 -2560
rect 1492 -2602 1532 -2562
rect 360 -2760 400 -2720
rect 1320 -2730 1360 -2690
rect -200 -3240 -160 -3200
<< metal1 >>
rect -320 510 -220 540
rect -320 470 -270 510
rect -230 470 -220 510
rect -320 440 -220 470
rect 430 510 890 540
rect 430 470 500 510
rect 540 470 600 510
rect 640 470 890 510
rect 430 440 890 470
rect 1530 510 1990 540
rect 1530 470 1560 510
rect 1600 470 1740 510
rect 1780 470 1920 510
rect 1960 470 1990 510
rect 1530 440 1990 470
rect 2630 500 2730 530
rect 2630 460 2660 500
rect 2700 460 2730 500
rect 2630 430 2730 460
rect -540 330 -460 360
rect -540 290 -520 330
rect -480 290 -460 330
rect -540 260 -460 290
rect 210 340 290 370
rect 210 300 230 340
rect 270 300 290 340
rect 210 270 290 300
rect 1310 340 1390 370
rect 1310 300 1330 340
rect 1370 300 1390 340
rect 530 260 610 280
rect 530 220 550 260
rect 590 220 610 260
rect 530 200 610 220
rect 890 260 970 290
rect 1310 270 1390 300
rect 2410 330 2490 360
rect 2410 290 2430 330
rect 2470 290 2490 330
rect 890 220 910 260
rect 950 220 970 260
rect 890 200 970 220
rect -220 180 -140 200
rect -220 140 -200 180
rect -160 140 -140 180
rect -220 100 -140 140
rect -220 60 -200 100
rect -160 60 -140 100
rect -220 -180 -140 60
rect 530 180 970 200
rect 530 140 550 180
rect 590 140 910 180
rect 950 140 970 180
rect 530 120 970 140
rect 530 100 610 120
rect 530 60 550 100
rect 590 60 610 100
rect 530 40 610 60
rect 890 100 970 120
rect 890 60 910 100
rect 950 60 970 100
rect 890 50 970 60
rect 1450 260 1530 280
rect 1450 220 1470 260
rect 1510 220 1530 260
rect 1450 200 1530 220
rect 1810 260 1890 280
rect 1810 220 1830 260
rect 1870 220 1890 260
rect 1810 200 1890 220
rect 1450 180 1890 200
rect 1450 140 1470 180
rect 1510 140 1830 180
rect 1870 140 1890 180
rect 1450 120 1890 140
rect 1450 100 1530 120
rect 1450 60 1470 100
rect 1510 60 1530 100
rect 1450 40 1530 60
rect 1810 100 1890 120
rect 1810 60 1830 100
rect 1870 60 1890 100
rect 1810 40 1890 60
rect 2410 -180 2490 290
rect 2550 170 2630 190
rect 2550 130 2570 170
rect 2610 130 2630 170
rect 2550 90 2630 130
rect 2550 50 2570 90
rect 2610 50 2630 90
rect 2550 -180 2630 50
rect -220 -280 2630 -180
rect -540 -770 -460 -740
rect -540 -810 -520 -770
rect -480 -810 -460 -770
rect -540 -840 -460 -810
rect 190 -760 1770 -660
rect 190 -1630 290 -760
rect 1490 -800 1770 -760
rect 1490 -840 1500 -800
rect 1540 -840 1720 -800
rect 1760 -840 1770 -800
rect 1490 -870 1770 -840
rect 2230 -870 2310 -770
rect 420 -970 500 -940
rect 420 -1010 440 -970
rect 480 -1010 500 -970
rect 420 -1040 500 -1010
rect 1270 -970 1350 -940
rect 1270 -1010 1290 -970
rect 1330 -1010 1350 -970
rect 1270 -1040 1350 -1010
rect 640 -1460 920 -1430
rect 640 -1500 710 -1460
rect 750 -1500 810 -1460
rect 850 -1500 920 -1460
rect 640 -1530 920 -1500
rect -320 -1660 290 -1630
rect -320 -1700 -310 -1660
rect -270 -1700 -90 -1660
rect -50 -1700 290 -1660
rect -320 -1730 290 -1700
rect 190 -2040 290 -1730
rect 740 -1660 820 -1530
rect 2450 -1660 2730 -1640
rect 740 -1670 2730 -1660
rect 740 -1710 2460 -1670
rect 2500 -1710 2680 -1670
rect 2720 -1710 2730 -1670
rect 740 -1740 2730 -1710
rect 190 -2140 1110 -2040
rect 340 -2380 420 -2350
rect 340 -2420 360 -2380
rect 400 -2420 420 -2380
rect 1030 -2410 1110 -2140
rect 340 -2450 420 -2420
rect 670 -2438 1110 -2410
rect 670 -2478 696 -2438
rect 736 -2478 1110 -2438
rect 1300 -2380 1380 -2350
rect 1300 -2420 1320 -2380
rect 1360 -2420 1380 -2380
rect 1300 -2450 1380 -2420
rect 1560 -2430 1640 -2390
rect 2050 -2430 2130 -1740
rect 1560 -2440 2130 -2430
rect 670 -2500 1110 -2478
rect 170 -2560 570 -2540
rect 170 -2600 520 -2560
rect 560 -2600 570 -2560
rect 170 -2620 570 -2600
rect 1030 -2550 1110 -2500
rect 1560 -2480 1580 -2440
rect 1620 -2480 2130 -2440
rect 1560 -2510 2130 -2480
rect 1030 -2562 1550 -2550
rect 1030 -2602 1492 -2562
rect 1532 -2602 1550 -2562
rect 1030 -2630 1550 -2602
rect 1300 -2690 1380 -2660
rect 340 -2720 420 -2690
rect 340 -2760 360 -2720
rect 400 -2760 420 -2720
rect 1300 -2730 1320 -2690
rect 1360 -2730 1380 -2690
rect 1300 -2760 1380 -2730
rect 340 -2790 420 -2760
rect -220 -3200 105 -3190
rect -220 -3240 -200 -3200
rect -160 -3240 105 -3200
rect -220 -3260 105 -3240
use sky130_fd_pr__res_xhigh_po_0p35_R469US  sky130_fd_pr__res_xhigh_po_0p35_R469US_0
timestamp 1726131431
transform 0 -1 1342 1 0 -3225
box -35 -1272 35 1272
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 478 0 1 -2822
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 1458 0 1 -2822
box -38 -48 314 592
<< labels >>
rlabel metal1 190 -2540 190 -2540 1 Dctrl
port 1 n
rlabel metal1 -260 540 -260 540 1 Vbs1
port 2 n
rlabel metal1 2680 530 2680 530 1 Vbs2
port 3 n
rlabel metal1 560 540 560 540 1 Vbs3
port 4 n
rlabel metal1 1760 540 1760 540 1 Vbs4
port 5 n
rlabel locali 3010 90 3010 90 1 Isup
port 6 n
rlabel locali -500 840 -500 840 1 VCCA
port 7 n
rlabel metal1 -70 -3230 -60 -3220 1 input_R
<< end >>
