magic
tech sky130A
timestamp 1726473936
<< nwell >>
rect -290 -40 -50 220
rect 85 -40 505 220
rect 635 -40 1055 220
rect 1185 -45 1425 215
rect -290 -815 40 -335
rect 1095 -820 1425 -340
<< pwell >>
rect 190 -715 520 -435
rect 630 -715 960 -435
<< nmos >>
rect 320 -675 370 -475
rect 410 -675 460 -475
rect 760 -675 810 -475
rect 850 -675 900 -475
<< pmoshvt >>
rect -160 0 -110 180
rect 215 0 265 180
rect 305 0 355 180
rect 395 0 445 180
rect 765 0 815 180
rect 855 0 905 180
rect 945 0 995 180
rect 1315 -5 1365 175
rect -160 -775 -110 -375
rect -70 -775 -20 -375
rect 1225 -780 1275 -380
rect 1315 -780 1365 -380
<< ndiff >>
rect 280 -490 320 -475
rect 280 -510 290 -490
rect 310 -510 320 -490
rect 280 -530 320 -510
rect 280 -550 290 -530
rect 310 -550 320 -530
rect 280 -570 320 -550
rect 280 -590 290 -570
rect 310 -590 320 -570
rect 280 -610 320 -590
rect 280 -630 290 -610
rect 310 -630 320 -610
rect 280 -675 320 -630
rect 370 -490 410 -475
rect 370 -510 380 -490
rect 400 -510 410 -490
rect 370 -530 410 -510
rect 370 -550 380 -530
rect 400 -550 410 -530
rect 370 -570 410 -550
rect 370 -590 380 -570
rect 400 -590 410 -570
rect 370 -610 410 -590
rect 370 -630 380 -610
rect 400 -630 410 -610
rect 370 -675 410 -630
rect 460 -490 500 -475
rect 460 -510 470 -490
rect 490 -510 500 -490
rect 460 -530 500 -510
rect 720 -490 760 -475
rect 720 -510 730 -490
rect 750 -510 760 -490
rect 460 -550 470 -530
rect 490 -550 500 -530
rect 460 -570 500 -550
rect 460 -590 470 -570
rect 490 -590 500 -570
rect 460 -610 500 -590
rect 460 -630 470 -610
rect 490 -630 500 -610
rect 460 -675 500 -630
rect 720 -530 760 -510
rect 720 -550 730 -530
rect 750 -550 760 -530
rect 720 -570 760 -550
rect 720 -590 730 -570
rect 750 -590 760 -570
rect 720 -610 760 -590
rect 720 -630 730 -610
rect 750 -630 760 -610
rect 720 -675 760 -630
rect 810 -490 850 -475
rect 810 -510 820 -490
rect 840 -510 850 -490
rect 810 -530 850 -510
rect 810 -550 820 -530
rect 840 -550 850 -530
rect 810 -570 850 -550
rect 810 -590 820 -570
rect 840 -590 850 -570
rect 810 -610 850 -590
rect 810 -630 820 -610
rect 840 -630 850 -610
rect 810 -675 850 -630
rect 900 -490 940 -475
rect 900 -510 910 -490
rect 930 -510 940 -490
rect 900 -530 940 -510
rect 900 -550 910 -530
rect 930 -550 940 -530
rect 900 -570 940 -550
rect 900 -590 910 -570
rect 930 -590 940 -570
rect 900 -610 940 -590
rect 900 -630 910 -610
rect 930 -630 940 -610
rect 900 -675 940 -630
<< pdiff >>
rect -200 170 -160 180
rect -200 150 -190 170
rect -170 150 -160 170
rect -200 130 -160 150
rect -200 110 -190 130
rect -170 110 -160 130
rect -200 90 -160 110
rect -200 70 -190 90
rect -170 70 -160 90
rect -200 50 -160 70
rect -200 30 -190 50
rect -170 30 -160 50
rect -200 0 -160 30
rect -110 170 -70 180
rect -110 150 -100 170
rect -80 150 -70 170
rect -110 130 -70 150
rect 175 170 215 180
rect 175 150 185 170
rect 205 150 215 170
rect -110 110 -100 130
rect -80 110 -70 130
rect -110 90 -70 110
rect -110 70 -100 90
rect -80 70 -70 90
rect -110 50 -70 70
rect -110 30 -100 50
rect -80 30 -70 50
rect -110 0 -70 30
rect 175 130 215 150
rect 175 110 185 130
rect 205 110 215 130
rect 175 90 215 110
rect 175 70 185 90
rect 205 70 215 90
rect 175 50 215 70
rect 175 30 185 50
rect 205 30 215 50
rect 175 0 215 30
rect 265 170 305 180
rect 265 150 275 170
rect 295 150 305 170
rect 265 130 305 150
rect 265 110 275 130
rect 295 110 305 130
rect 265 90 305 110
rect 265 70 275 90
rect 295 70 305 90
rect 265 50 305 70
rect 265 30 275 50
rect 295 30 305 50
rect 265 0 305 30
rect 355 170 395 180
rect 355 150 365 170
rect 385 150 395 170
rect 355 130 395 150
rect 355 110 365 130
rect 385 110 395 130
rect 355 90 395 110
rect 355 70 365 90
rect 385 70 395 90
rect 355 50 395 70
rect 355 30 365 50
rect 385 30 395 50
rect 355 0 395 30
rect 445 170 485 180
rect 445 150 455 170
rect 475 150 485 170
rect 445 130 485 150
rect 725 170 765 180
rect 725 150 735 170
rect 755 150 765 170
rect 445 110 455 130
rect 475 110 485 130
rect 445 90 485 110
rect 445 70 455 90
rect 475 70 485 90
rect 445 50 485 70
rect 445 30 455 50
rect 475 30 485 50
rect 445 0 485 30
rect 725 130 765 150
rect 725 110 735 130
rect 755 110 765 130
rect 725 90 765 110
rect 725 70 735 90
rect 755 70 765 90
rect 725 50 765 70
rect 725 30 735 50
rect 755 30 765 50
rect 725 0 765 30
rect 815 170 855 180
rect 815 150 825 170
rect 845 150 855 170
rect 815 130 855 150
rect 815 110 825 130
rect 845 110 855 130
rect 815 90 855 110
rect 815 70 825 90
rect 845 70 855 90
rect 815 50 855 70
rect 815 30 825 50
rect 845 30 855 50
rect 815 0 855 30
rect 905 170 945 180
rect 905 150 915 170
rect 935 150 945 170
rect 905 130 945 150
rect 905 110 915 130
rect 935 110 945 130
rect 905 90 945 110
rect 905 70 915 90
rect 935 70 945 90
rect 905 50 945 70
rect 905 30 915 50
rect 935 30 945 50
rect 905 0 945 30
rect 995 170 1035 180
rect 995 150 1005 170
rect 1025 150 1035 170
rect 995 130 1035 150
rect 1275 165 1315 175
rect 1275 145 1285 165
rect 1305 145 1315 165
rect 995 110 1005 130
rect 1025 110 1035 130
rect 995 90 1035 110
rect 995 70 1005 90
rect 1025 70 1035 90
rect 995 50 1035 70
rect 995 30 1005 50
rect 1025 30 1035 50
rect 995 0 1035 30
rect 1275 125 1315 145
rect 1275 105 1285 125
rect 1305 105 1315 125
rect 1275 85 1315 105
rect 1275 65 1285 85
rect 1305 65 1315 85
rect 1275 45 1315 65
rect 1275 25 1285 45
rect 1305 25 1315 45
rect 1275 -5 1315 25
rect 1365 165 1405 175
rect 1365 145 1375 165
rect 1395 145 1405 165
rect 1365 125 1405 145
rect 1365 105 1375 125
rect 1395 105 1405 125
rect 1365 85 1405 105
rect 1365 65 1375 85
rect 1395 65 1405 85
rect 1365 45 1405 65
rect 1365 25 1375 45
rect 1395 25 1405 45
rect 1365 -5 1405 25
rect -200 -385 -160 -375
rect -200 -405 -190 -385
rect -170 -405 -160 -385
rect -200 -425 -160 -405
rect -200 -445 -190 -425
rect -170 -445 -160 -425
rect -200 -465 -160 -445
rect -200 -485 -190 -465
rect -170 -485 -160 -465
rect -200 -505 -160 -485
rect -200 -525 -190 -505
rect -170 -525 -160 -505
rect -200 -545 -160 -525
rect -200 -565 -190 -545
rect -170 -565 -160 -545
rect -200 -585 -160 -565
rect -200 -605 -190 -585
rect -170 -605 -160 -585
rect -200 -625 -160 -605
rect -200 -645 -190 -625
rect -170 -645 -160 -625
rect -200 -665 -160 -645
rect -200 -685 -190 -665
rect -170 -685 -160 -665
rect -200 -705 -160 -685
rect -200 -725 -190 -705
rect -170 -725 -160 -705
rect -200 -745 -160 -725
rect -200 -765 -190 -745
rect -170 -765 -160 -745
rect -200 -775 -160 -765
rect -110 -385 -70 -375
rect -110 -405 -100 -385
rect -80 -405 -70 -385
rect -110 -425 -70 -405
rect -110 -445 -100 -425
rect -80 -445 -70 -425
rect -110 -465 -70 -445
rect -110 -485 -100 -465
rect -80 -485 -70 -465
rect -110 -505 -70 -485
rect -110 -525 -100 -505
rect -80 -525 -70 -505
rect -110 -545 -70 -525
rect -110 -565 -100 -545
rect -80 -565 -70 -545
rect -110 -585 -70 -565
rect -110 -605 -100 -585
rect -80 -605 -70 -585
rect -110 -625 -70 -605
rect -110 -645 -100 -625
rect -80 -645 -70 -625
rect -110 -665 -70 -645
rect -110 -685 -100 -665
rect -80 -685 -70 -665
rect -110 -705 -70 -685
rect -110 -725 -100 -705
rect -80 -725 -70 -705
rect -110 -745 -70 -725
rect -110 -765 -100 -745
rect -80 -765 -70 -745
rect -110 -775 -70 -765
rect -20 -385 20 -375
rect -20 -405 -10 -385
rect 10 -405 20 -385
rect -20 -425 20 -405
rect -20 -445 -10 -425
rect 10 -445 20 -425
rect 1185 -390 1225 -380
rect 1185 -410 1195 -390
rect 1215 -410 1225 -390
rect 1185 -430 1225 -410
rect -20 -465 20 -445
rect -20 -485 -10 -465
rect 10 -485 20 -465
rect -20 -505 20 -485
rect -20 -525 -10 -505
rect 10 -525 20 -505
rect -20 -545 20 -525
rect -20 -565 -10 -545
rect 10 -565 20 -545
rect -20 -585 20 -565
rect -20 -605 -10 -585
rect 10 -605 20 -585
rect -20 -625 20 -605
rect -20 -645 -10 -625
rect 10 -645 20 -625
rect -20 -665 20 -645
rect -20 -685 -10 -665
rect 10 -685 20 -665
rect 1185 -450 1195 -430
rect 1215 -450 1225 -430
rect 1185 -470 1225 -450
rect 1185 -490 1195 -470
rect 1215 -490 1225 -470
rect 1185 -510 1225 -490
rect 1185 -530 1195 -510
rect 1215 -530 1225 -510
rect 1185 -550 1225 -530
rect 1185 -570 1195 -550
rect 1215 -570 1225 -550
rect 1185 -590 1225 -570
rect 1185 -610 1195 -590
rect 1215 -610 1225 -590
rect 1185 -630 1225 -610
rect 1185 -650 1195 -630
rect 1215 -650 1225 -630
rect 1185 -670 1225 -650
rect -20 -705 20 -685
rect -20 -725 -10 -705
rect 10 -725 20 -705
rect -20 -745 20 -725
rect -20 -765 -10 -745
rect 10 -765 20 -745
rect 1185 -690 1195 -670
rect 1215 -690 1225 -670
rect 1185 -710 1225 -690
rect 1185 -730 1195 -710
rect 1215 -730 1225 -710
rect 1185 -750 1225 -730
rect -20 -775 20 -765
rect 1185 -770 1195 -750
rect 1215 -770 1225 -750
rect 1185 -780 1225 -770
rect 1275 -390 1315 -380
rect 1275 -410 1285 -390
rect 1305 -410 1315 -390
rect 1275 -430 1315 -410
rect 1275 -450 1285 -430
rect 1305 -450 1315 -430
rect 1275 -470 1315 -450
rect 1275 -490 1285 -470
rect 1305 -490 1315 -470
rect 1275 -510 1315 -490
rect 1275 -530 1285 -510
rect 1305 -530 1315 -510
rect 1275 -550 1315 -530
rect 1275 -570 1285 -550
rect 1305 -570 1315 -550
rect 1275 -590 1315 -570
rect 1275 -610 1285 -590
rect 1305 -610 1315 -590
rect 1275 -630 1315 -610
rect 1275 -650 1285 -630
rect 1305 -650 1315 -630
rect 1275 -670 1315 -650
rect 1275 -690 1285 -670
rect 1305 -690 1315 -670
rect 1275 -710 1315 -690
rect 1275 -730 1285 -710
rect 1305 -730 1315 -710
rect 1275 -750 1315 -730
rect 1275 -770 1285 -750
rect 1305 -770 1315 -750
rect 1275 -780 1315 -770
rect 1365 -390 1405 -380
rect 1365 -410 1375 -390
rect 1395 -410 1405 -390
rect 1365 -430 1405 -410
rect 1365 -450 1375 -430
rect 1395 -450 1405 -430
rect 1365 -470 1405 -450
rect 1365 -490 1375 -470
rect 1395 -490 1405 -470
rect 1365 -510 1405 -490
rect 1365 -530 1375 -510
rect 1395 -530 1405 -510
rect 1365 -550 1405 -530
rect 1365 -570 1375 -550
rect 1395 -570 1405 -550
rect 1365 -590 1405 -570
rect 1365 -610 1375 -590
rect 1395 -610 1405 -590
rect 1365 -630 1405 -610
rect 1365 -650 1375 -630
rect 1395 -650 1405 -630
rect 1365 -670 1405 -650
rect 1365 -690 1375 -670
rect 1395 -690 1405 -670
rect 1365 -710 1405 -690
rect 1365 -730 1375 -710
rect 1395 -730 1405 -710
rect 1365 -750 1405 -730
rect 1365 -770 1375 -750
rect 1395 -770 1405 -750
rect 1365 -780 1405 -770
<< ndiffc >>
rect 290 -510 310 -490
rect 290 -550 310 -530
rect 290 -590 310 -570
rect 290 -630 310 -610
rect 380 -510 400 -490
rect 380 -550 400 -530
rect 380 -590 400 -570
rect 380 -630 400 -610
rect 470 -510 490 -490
rect 730 -510 750 -490
rect 470 -550 490 -530
rect 470 -590 490 -570
rect 470 -630 490 -610
rect 730 -550 750 -530
rect 730 -590 750 -570
rect 730 -630 750 -610
rect 820 -510 840 -490
rect 820 -550 840 -530
rect 820 -590 840 -570
rect 820 -630 840 -610
rect 910 -510 930 -490
rect 910 -550 930 -530
rect 910 -590 930 -570
rect 910 -630 930 -610
<< pdiffc >>
rect -190 150 -170 170
rect -190 110 -170 130
rect -190 70 -170 90
rect -190 30 -170 50
rect -100 150 -80 170
rect 185 150 205 170
rect -100 110 -80 130
rect -100 70 -80 90
rect -100 30 -80 50
rect 185 110 205 130
rect 185 70 205 90
rect 185 30 205 50
rect 275 150 295 170
rect 275 110 295 130
rect 275 70 295 90
rect 275 30 295 50
rect 365 150 385 170
rect 365 110 385 130
rect 365 70 385 90
rect 365 30 385 50
rect 455 150 475 170
rect 735 150 755 170
rect 455 110 475 130
rect 455 70 475 90
rect 455 30 475 50
rect 735 110 755 130
rect 735 70 755 90
rect 735 30 755 50
rect 825 150 845 170
rect 825 110 845 130
rect 825 70 845 90
rect 825 30 845 50
rect 915 150 935 170
rect 915 110 935 130
rect 915 70 935 90
rect 915 30 935 50
rect 1005 150 1025 170
rect 1285 145 1305 165
rect 1005 110 1025 130
rect 1005 70 1025 90
rect 1005 30 1025 50
rect 1285 105 1305 125
rect 1285 65 1305 85
rect 1285 25 1305 45
rect 1375 145 1395 165
rect 1375 105 1395 125
rect 1375 65 1395 85
rect 1375 25 1395 45
rect -190 -405 -170 -385
rect -190 -445 -170 -425
rect -190 -485 -170 -465
rect -190 -525 -170 -505
rect -190 -565 -170 -545
rect -190 -605 -170 -585
rect -190 -645 -170 -625
rect -190 -685 -170 -665
rect -190 -725 -170 -705
rect -190 -765 -170 -745
rect -100 -405 -80 -385
rect -100 -445 -80 -425
rect -100 -485 -80 -465
rect -100 -525 -80 -505
rect -100 -565 -80 -545
rect -100 -605 -80 -585
rect -100 -645 -80 -625
rect -100 -685 -80 -665
rect -100 -725 -80 -705
rect -100 -765 -80 -745
rect -10 -405 10 -385
rect -10 -445 10 -425
rect 1195 -410 1215 -390
rect -10 -485 10 -465
rect -10 -525 10 -505
rect -10 -565 10 -545
rect -10 -605 10 -585
rect -10 -645 10 -625
rect -10 -685 10 -665
rect 1195 -450 1215 -430
rect 1195 -490 1215 -470
rect 1195 -530 1215 -510
rect 1195 -570 1215 -550
rect 1195 -610 1215 -590
rect 1195 -650 1215 -630
rect -10 -725 10 -705
rect -10 -765 10 -745
rect 1195 -690 1215 -670
rect 1195 -730 1215 -710
rect 1195 -770 1215 -750
rect 1285 -410 1305 -390
rect 1285 -450 1305 -430
rect 1285 -490 1305 -470
rect 1285 -530 1305 -510
rect 1285 -570 1305 -550
rect 1285 -610 1305 -590
rect 1285 -650 1305 -630
rect 1285 -690 1305 -670
rect 1285 -730 1305 -710
rect 1285 -770 1305 -750
rect 1375 -410 1395 -390
rect 1375 -450 1395 -430
rect 1375 -490 1395 -470
rect 1375 -530 1395 -510
rect 1375 -570 1395 -550
rect 1375 -610 1395 -590
rect 1375 -650 1395 -630
rect 1375 -690 1395 -670
rect 1375 -730 1395 -710
rect 1375 -770 1395 -750
<< psubdiff >>
rect 210 -485 250 -470
rect 210 -505 220 -485
rect 240 -505 250 -485
rect 210 -520 250 -505
rect 650 -485 690 -470
rect 650 -505 660 -485
rect 680 -505 690 -485
rect 650 -520 690 -505
<< nsubdiff >>
rect -270 165 -230 180
rect -270 145 -260 165
rect -240 145 -230 165
rect -270 130 -230 145
rect 105 170 145 185
rect 105 150 115 170
rect 135 150 145 170
rect 105 135 145 150
rect 655 170 695 185
rect 655 150 665 170
rect 685 150 695 170
rect 655 135 695 150
rect 1205 165 1245 180
rect 1205 145 1215 165
rect 1235 145 1245 165
rect 1205 130 1245 145
rect -270 -385 -230 -370
rect -270 -405 -260 -385
rect -240 -405 -230 -385
rect -270 -420 -230 -405
rect 1115 -400 1155 -385
rect 1115 -420 1125 -400
rect 1145 -420 1155 -400
rect 1115 -435 1155 -420
<< psubdiffcont >>
rect 220 -505 240 -485
rect 660 -505 680 -485
<< nsubdiffcont >>
rect -260 145 -240 165
rect 115 150 135 170
rect 665 150 685 170
rect 1215 145 1235 165
rect -260 -405 -240 -385
rect 1125 -420 1145 -400
<< poly >>
rect -160 255 -110 270
rect -160 235 -135 255
rect -115 235 -110 255
rect -160 180 -110 235
rect 215 255 445 270
rect 215 235 250 255
rect 270 235 300 255
rect 320 235 445 255
rect 215 220 445 235
rect 215 180 265 220
rect 305 180 355 220
rect 395 180 445 220
rect 765 255 995 270
rect 765 235 780 255
rect 800 235 870 255
rect 890 235 960 255
rect 980 235 995 255
rect 765 220 995 235
rect 765 180 815 220
rect 855 180 905 220
rect 945 180 995 220
rect 1315 250 1365 265
rect 1315 230 1330 250
rect 1350 230 1365 250
rect 1315 175 1365 230
rect -160 -40 -110 0
rect 215 -40 265 0
rect 305 -40 355 0
rect 395 -40 445 0
rect 765 -40 815 0
rect 855 -40 905 0
rect 945 -40 995 0
rect 1315 -45 1365 -5
rect -160 -375 -110 -335
rect -70 -375 -20 -335
rect 1225 -380 1275 -340
rect 1315 -380 1365 -340
rect 760 -400 900 -385
rect 760 -420 795 -400
rect 815 -420 840 -400
rect 860 -420 900 -400
rect 760 -435 900 -420
rect 320 -475 370 -435
rect 410 -475 460 -435
rect 760 -475 810 -435
rect 850 -475 900 -435
rect 320 -715 370 -675
rect 410 -715 460 -675
rect 760 -715 810 -675
rect 850 -715 900 -675
rect 320 -730 460 -715
rect 320 -750 355 -730
rect 375 -750 405 -730
rect 425 -750 460 -730
rect 320 -765 460 -750
rect -160 -815 -110 -775
rect -70 -815 -20 -775
rect -160 -830 -20 -815
rect -160 -850 -155 -830
rect -135 -850 -45 -830
rect -25 -850 -20 -830
rect -160 -865 -20 -850
rect 1225 -820 1275 -780
rect 1315 -820 1365 -780
rect 1225 -835 1365 -820
rect 1225 -855 1230 -835
rect 1250 -855 1340 -835
rect 1360 -855 1365 -835
rect 1225 -870 1365 -855
<< polycont >>
rect -135 235 -115 255
rect 250 235 270 255
rect 300 235 320 255
rect 780 235 800 255
rect 870 235 890 255
rect 960 235 980 255
rect 1330 230 1350 250
rect 795 -420 815 -400
rect 840 -420 860 -400
rect 355 -750 375 -730
rect 405 -750 425 -730
rect -155 -850 -135 -830
rect -45 -850 -25 -830
rect 1230 -855 1250 -835
rect 1340 -855 1360 -835
<< locali >>
rect -270 165 -230 370
rect -270 145 -260 165
rect -240 145 -230 165
rect -270 130 -230 145
rect -200 170 -160 370
rect -140 255 -110 270
rect -140 235 -135 255
rect -115 235 -110 255
rect -140 220 -110 235
rect -200 150 -190 170
rect -170 150 -160 170
rect -200 130 -160 150
rect -200 110 -190 130
rect -170 110 -160 130
rect -200 90 -160 110
rect -200 70 -190 90
rect -170 70 -160 90
rect -200 50 -160 70
rect -200 30 -190 50
rect -170 30 -160 50
rect -200 0 -160 30
rect -110 170 -70 180
rect -110 150 -100 170
rect -80 150 -70 170
rect -110 130 -70 150
rect 105 170 145 370
rect 105 150 115 170
rect 135 150 145 170
rect 105 135 145 150
rect 175 330 395 370
rect 175 170 215 330
rect 235 255 335 270
rect 235 235 250 255
rect 270 235 300 255
rect 320 235 335 255
rect 235 220 335 235
rect 175 150 185 170
rect 205 150 215 170
rect -110 110 -100 130
rect -80 110 -70 130
rect -110 90 -70 110
rect -110 70 -100 90
rect -80 70 -70 90
rect -110 50 -70 70
rect -110 30 -100 50
rect -80 30 -70 50
rect -110 0 -70 30
rect 175 130 215 150
rect 175 110 185 130
rect 205 110 215 130
rect 175 90 215 110
rect 175 70 185 90
rect 205 70 215 90
rect 175 50 215 70
rect 175 30 185 50
rect 205 30 215 50
rect 175 0 215 30
rect 265 170 305 180
rect 265 150 275 170
rect 295 150 305 170
rect 265 130 305 150
rect 265 110 275 130
rect 295 110 305 130
rect 265 90 305 110
rect 265 70 275 90
rect 295 70 305 90
rect 265 50 305 70
rect 265 30 275 50
rect 295 30 305 50
rect 265 0 305 30
rect 355 170 395 330
rect 765 255 995 270
rect 765 235 780 255
rect 800 235 870 255
rect 890 235 960 255
rect 980 235 995 255
rect 765 220 995 235
rect 1315 250 1365 265
rect 1315 230 1330 250
rect 1350 230 1365 250
rect 1315 215 1365 230
rect 355 150 365 170
rect 385 150 395 170
rect 355 130 395 150
rect 355 110 365 130
rect 385 110 395 130
rect 355 90 395 110
rect 355 70 365 90
rect 385 70 395 90
rect 355 50 395 70
rect 355 30 365 50
rect 385 30 395 50
rect 355 0 395 30
rect 445 170 485 180
rect 445 150 455 170
rect 475 150 485 170
rect 445 130 485 150
rect 445 110 455 130
rect 475 110 485 130
rect 445 90 485 110
rect 655 170 695 185
rect 655 150 665 170
rect 685 150 695 170
rect 655 100 695 150
rect 725 170 765 180
rect 725 150 735 170
rect 755 150 765 170
rect 725 130 765 150
rect 725 110 735 130
rect 755 110 765 130
rect 445 70 455 90
rect 475 70 485 90
rect 445 50 485 70
rect 445 30 455 50
rect 475 30 485 50
rect 445 0 485 30
rect 725 90 765 110
rect 725 70 735 90
rect 755 70 765 90
rect 725 50 765 70
rect 725 30 735 50
rect 755 30 765 50
rect 725 0 765 30
rect 815 170 855 180
rect 815 150 825 170
rect 845 150 855 170
rect 815 130 855 150
rect 815 110 825 130
rect 845 110 855 130
rect 815 90 855 110
rect 815 70 825 90
rect 845 70 855 90
rect 815 50 855 70
rect 815 30 825 50
rect 845 30 855 50
rect 815 -75 855 30
rect 905 170 945 180
rect 905 150 915 170
rect 935 150 945 170
rect 905 130 945 150
rect 905 110 915 130
rect 935 110 945 130
rect 905 90 945 110
rect 905 70 915 90
rect 935 70 945 90
rect 905 50 945 70
rect 905 30 915 50
rect 935 30 945 50
rect 905 0 945 30
rect 995 170 1035 180
rect 995 150 1005 170
rect 1025 150 1035 170
rect 995 130 1035 150
rect 1205 165 1245 180
rect 1205 145 1215 165
rect 1235 145 1245 165
rect 1205 130 1245 145
rect 1275 165 1315 175
rect 1275 145 1285 165
rect 1305 145 1315 165
rect 995 110 1005 130
rect 1025 110 1035 130
rect 995 90 1035 110
rect 995 70 1005 90
rect 1025 70 1035 90
rect 995 50 1035 70
rect 995 30 1005 50
rect 1025 30 1035 50
rect 995 -75 1035 30
rect 1275 125 1315 145
rect 1275 105 1285 125
rect 1305 105 1315 125
rect 1275 85 1315 105
rect 1275 65 1285 85
rect 1305 65 1315 85
rect 1275 45 1315 65
rect 1275 25 1285 45
rect 1305 25 1315 45
rect 1275 -5 1315 25
rect 1365 165 1405 175
rect 1365 145 1375 165
rect 1395 145 1405 165
rect 1365 125 1405 145
rect 1365 105 1375 125
rect 1395 105 1405 125
rect 1365 85 1405 105
rect 1365 65 1375 85
rect 1395 65 1405 85
rect 1365 45 1405 65
rect 1365 25 1375 45
rect 1395 25 1475 45
rect 1365 -5 1475 25
rect 815 -115 1035 -75
rect -200 -270 20 -230
rect 720 -270 940 -230
rect 1185 -270 1405 -230
rect -270 -385 -230 -270
rect -270 -405 -260 -385
rect -240 -405 -230 -385
rect -270 -420 -230 -405
rect -200 -385 -160 -270
rect -200 -405 -190 -385
rect -170 -405 -160 -385
rect -200 -425 -160 -405
rect -200 -445 -190 -425
rect -170 -445 -160 -425
rect -200 -465 -160 -445
rect -200 -485 -190 -465
rect -170 -485 -160 -465
rect -200 -505 -160 -485
rect -200 -525 -190 -505
rect -170 -525 -160 -505
rect -200 -545 -160 -525
rect -200 -565 -190 -545
rect -170 -565 -160 -545
rect -200 -585 -160 -565
rect -200 -605 -190 -585
rect -170 -605 -160 -585
rect -200 -625 -160 -605
rect -200 -645 -190 -625
rect -170 -645 -160 -625
rect -200 -665 -160 -645
rect -200 -685 -190 -665
rect -170 -685 -160 -665
rect -200 -705 -160 -685
rect -200 -725 -190 -705
rect -170 -725 -160 -705
rect -200 -745 -160 -725
rect -200 -765 -190 -745
rect -170 -765 -160 -745
rect -200 -775 -160 -765
rect -110 -385 -70 -375
rect -110 -405 -100 -385
rect -80 -405 -70 -385
rect -110 -425 -70 -405
rect -110 -445 -100 -425
rect -80 -445 -70 -425
rect -110 -465 -70 -445
rect -110 -485 -100 -465
rect -80 -485 -70 -465
rect -110 -505 -70 -485
rect -110 -525 -100 -505
rect -80 -525 -70 -505
rect -110 -545 -70 -525
rect -110 -565 -100 -545
rect -80 -565 -70 -545
rect -110 -585 -70 -565
rect -110 -605 -100 -585
rect -80 -605 -70 -585
rect -110 -625 -70 -605
rect -110 -645 -100 -625
rect -80 -645 -70 -625
rect -110 -665 -70 -645
rect -110 -685 -100 -665
rect -80 -685 -70 -665
rect -110 -705 -70 -685
rect -110 -725 -100 -705
rect -80 -725 -70 -705
rect -110 -745 -70 -725
rect -110 -765 -100 -745
rect -80 -765 -70 -745
rect -110 -775 -70 -765
rect -20 -385 20 -270
rect -20 -405 -10 -385
rect 10 -405 20 -385
rect -20 -425 20 -405
rect -20 -445 -10 -425
rect 10 -445 20 -425
rect -20 -465 20 -445
rect -20 -485 -10 -465
rect 10 -485 20 -465
rect -20 -505 20 -485
rect -20 -525 -10 -505
rect 10 -525 20 -505
rect -20 -545 20 -525
rect -20 -565 -10 -545
rect 10 -565 20 -545
rect -20 -585 20 -565
rect -20 -605 -10 -585
rect 10 -605 20 -585
rect -20 -625 20 -605
rect -20 -645 -10 -625
rect 10 -645 20 -625
rect -20 -665 20 -645
rect -20 -685 -10 -665
rect 10 -685 20 -665
rect -20 -705 20 -685
rect -20 -725 -10 -705
rect 10 -725 20 -705
rect -20 -745 20 -725
rect -20 -765 -10 -745
rect 10 -765 20 -745
rect -20 -775 20 -765
rect 210 -485 250 -470
rect 210 -505 220 -485
rect 240 -505 250 -485
rect -160 -830 -130 -815
rect -160 -850 -155 -830
rect -135 -850 -130 -830
rect -160 -865 -130 -850
rect -50 -830 -20 -815
rect -50 -850 -45 -830
rect -25 -850 -20 -830
rect -50 -865 -20 -850
rect 210 -915 250 -505
rect 280 -490 320 -475
rect 280 -510 290 -490
rect 310 -510 320 -490
rect 280 -530 320 -510
rect 280 -550 290 -530
rect 310 -550 320 -530
rect 280 -570 320 -550
rect 280 -590 290 -570
rect 310 -590 320 -570
rect 280 -610 320 -590
rect 280 -630 290 -610
rect 310 -630 320 -610
rect 280 -875 320 -630
rect 370 -490 410 -270
rect 370 -510 380 -490
rect 400 -510 410 -490
rect 370 -530 410 -510
rect 370 -550 380 -530
rect 400 -550 410 -530
rect 370 -570 410 -550
rect 370 -590 380 -570
rect 400 -590 410 -570
rect 370 -610 410 -590
rect 370 -630 380 -610
rect 400 -630 410 -610
rect 370 -675 410 -630
rect 460 -490 500 -475
rect 460 -510 470 -490
rect 490 -510 500 -490
rect 460 -530 500 -510
rect 650 -485 690 -385
rect 650 -505 660 -485
rect 680 -505 690 -485
rect 650 -520 690 -505
rect 720 -490 760 -270
rect 785 -400 870 -385
rect 785 -420 795 -400
rect 815 -420 840 -400
rect 860 -420 870 -400
rect 785 -435 870 -420
rect 720 -510 730 -490
rect 750 -510 760 -490
rect 460 -550 470 -530
rect 490 -550 500 -530
rect 460 -570 500 -550
rect 460 -590 470 -570
rect 490 -590 500 -570
rect 460 -610 500 -590
rect 460 -630 470 -610
rect 490 -630 500 -610
rect 340 -730 440 -715
rect 340 -750 355 -730
rect 375 -750 405 -730
rect 425 -750 440 -730
rect 340 -765 440 -750
rect 460 -875 500 -630
rect 720 -530 760 -510
rect 720 -550 730 -530
rect 750 -550 760 -530
rect 720 -570 760 -550
rect 720 -590 730 -570
rect 750 -590 760 -570
rect 720 -610 760 -590
rect 720 -630 730 -610
rect 750 -630 760 -610
rect 720 -675 760 -630
rect 810 -490 850 -475
rect 810 -510 820 -490
rect 840 -510 850 -490
rect 810 -530 850 -510
rect 810 -550 820 -530
rect 840 -550 850 -530
rect 810 -570 850 -550
rect 810 -590 820 -570
rect 840 -590 850 -570
rect 810 -610 850 -590
rect 810 -630 820 -610
rect 840 -630 850 -610
rect 810 -850 850 -630
rect 900 -490 940 -270
rect 1115 -400 1155 -270
rect 1115 -420 1125 -400
rect 1145 -420 1155 -400
rect 1115 -435 1155 -420
rect 1185 -390 1225 -270
rect 1185 -410 1195 -390
rect 1215 -410 1225 -390
rect 1185 -430 1225 -410
rect 900 -510 910 -490
rect 930 -510 940 -490
rect 900 -530 940 -510
rect 900 -550 910 -530
rect 930 -550 940 -530
rect 900 -570 940 -550
rect 900 -590 910 -570
rect 930 -590 940 -570
rect 900 -610 940 -590
rect 900 -630 910 -610
rect 930 -630 940 -610
rect 900 -675 940 -630
rect 1185 -450 1195 -430
rect 1215 -450 1225 -430
rect 1185 -470 1225 -450
rect 1185 -490 1195 -470
rect 1215 -490 1225 -470
rect 1185 -510 1225 -490
rect 1185 -530 1195 -510
rect 1215 -530 1225 -510
rect 1185 -550 1225 -530
rect 1185 -570 1195 -550
rect 1215 -570 1225 -550
rect 1185 -590 1225 -570
rect 1185 -610 1195 -590
rect 1215 -610 1225 -590
rect 1185 -630 1225 -610
rect 1185 -650 1195 -630
rect 1215 -650 1225 -630
rect 1185 -670 1225 -650
rect 1185 -690 1195 -670
rect 1215 -690 1225 -670
rect 1185 -710 1225 -690
rect 1185 -730 1195 -710
rect 1215 -730 1225 -710
rect 1185 -750 1225 -730
rect 1185 -770 1195 -750
rect 1215 -770 1225 -750
rect 1185 -780 1225 -770
rect 1275 -390 1315 -380
rect 1275 -410 1285 -390
rect 1305 -410 1315 -390
rect 1275 -430 1315 -410
rect 1275 -450 1285 -430
rect 1305 -450 1315 -430
rect 1275 -470 1315 -450
rect 1275 -490 1285 -470
rect 1305 -490 1315 -470
rect 1275 -510 1315 -490
rect 1275 -530 1285 -510
rect 1305 -530 1315 -510
rect 1275 -550 1315 -530
rect 1275 -570 1285 -550
rect 1305 -570 1315 -550
rect 1275 -590 1315 -570
rect 1275 -610 1285 -590
rect 1305 -610 1315 -590
rect 1275 -630 1315 -610
rect 1275 -650 1285 -630
rect 1305 -650 1315 -630
rect 1275 -670 1315 -650
rect 1275 -690 1285 -670
rect 1305 -690 1315 -670
rect 1275 -710 1315 -690
rect 1275 -730 1285 -710
rect 1305 -730 1315 -710
rect 1275 -750 1315 -730
rect 1275 -770 1285 -750
rect 1305 -770 1315 -750
rect 1225 -835 1255 -820
rect 1225 -855 1230 -835
rect 1250 -855 1255 -835
rect 1225 -870 1255 -855
rect 280 -915 500 -875
rect 1275 -915 1315 -770
rect 1365 -390 1405 -270
rect 1365 -410 1375 -390
rect 1395 -410 1405 -390
rect 1365 -430 1405 -410
rect 1365 -450 1375 -430
rect 1395 -450 1405 -430
rect 1365 -470 1405 -450
rect 1365 -490 1375 -470
rect 1395 -490 1405 -470
rect 1365 -510 1405 -490
rect 1365 -530 1375 -510
rect 1395 -530 1405 -510
rect 1365 -550 1405 -530
rect 1365 -570 1375 -550
rect 1395 -570 1405 -550
rect 1365 -590 1405 -570
rect 1365 -610 1375 -590
rect 1395 -610 1405 -590
rect 1365 -630 1405 -610
rect 1365 -650 1375 -630
rect 1395 -650 1405 -630
rect 1365 -670 1405 -650
rect 1365 -690 1375 -670
rect 1395 -690 1405 -670
rect 1365 -710 1405 -690
rect 1365 -730 1375 -710
rect 1395 -730 1405 -710
rect 1365 -750 1405 -730
rect 1365 -770 1375 -750
rect 1395 -770 1405 -750
rect 1365 -780 1405 -770
rect 1335 -835 1365 -820
rect 1335 -855 1340 -835
rect 1360 -855 1365 -835
rect 1335 -870 1365 -855
<< viali >>
rect -260 145 -240 165
rect -135 235 -115 255
rect 115 150 135 170
rect 250 235 270 255
rect 300 235 320 255
rect -100 70 -80 90
rect -100 30 -80 50
rect 275 110 295 130
rect 275 70 295 90
rect 275 30 295 50
rect 780 235 800 255
rect 870 235 890 255
rect 960 235 980 255
rect 1330 230 1350 250
rect 455 110 475 130
rect 665 150 685 170
rect 735 110 755 130
rect 455 70 475 90
rect 455 30 475 50
rect 735 70 755 90
rect 735 30 755 50
rect 915 110 935 130
rect 915 70 935 90
rect 915 30 935 50
rect 1215 145 1235 165
rect 1285 65 1305 85
rect 1285 25 1305 45
rect -260 -405 -240 -385
rect 220 -505 240 -485
rect -155 -850 -135 -830
rect -45 -850 -25 -830
rect 660 -505 680 -485
rect 795 -420 815 -400
rect 840 -420 860 -400
rect 355 -750 375 -730
rect 405 -750 425 -730
rect 1125 -420 1145 -400
rect 1230 -855 1250 -835
rect 1340 -855 1360 -835
<< metal1 >>
rect -160 255 -110 270
rect -160 235 -135 255
rect -115 235 -110 255
rect -160 220 -110 235
rect 215 255 445 270
rect 215 235 250 255
rect 270 235 300 255
rect 320 235 445 255
rect 215 220 445 235
rect 765 255 995 270
rect 765 235 780 255
rect 800 235 870 255
rect 890 235 960 255
rect 980 235 995 255
rect 765 220 995 235
rect 1315 250 1365 265
rect 1315 230 1330 250
rect 1350 230 1365 250
rect 1315 215 1365 230
rect -270 165 -230 180
rect -270 145 -260 165
rect -240 145 -230 165
rect -270 130 -230 145
rect 105 170 145 185
rect 105 150 115 170
rect 135 150 145 170
rect 105 135 145 150
rect 655 170 695 185
rect 655 150 665 170
rect 685 150 695 170
rect 265 130 305 140
rect 265 110 275 130
rect 295 110 305 130
rect 265 100 305 110
rect 445 130 485 145
rect 655 135 695 150
rect 1205 165 1245 180
rect 1205 145 1215 165
rect 1235 145 1245 165
rect 445 110 455 130
rect 475 110 485 130
rect 445 100 485 110
rect -110 90 -70 100
rect -110 70 -100 90
rect -80 70 -70 90
rect -110 50 -70 70
rect -110 30 -100 50
rect -80 30 -70 50
rect -110 -90 -70 30
rect 265 90 485 100
rect 265 70 275 90
rect 295 70 455 90
rect 475 70 485 90
rect 265 60 485 70
rect 265 50 305 60
rect 265 30 275 50
rect 295 30 305 50
rect 265 20 305 30
rect 445 50 485 60
rect 445 30 455 50
rect 475 30 485 50
rect 445 25 485 30
rect 725 130 765 140
rect 725 110 735 130
rect 755 110 765 130
rect 725 100 765 110
rect 905 130 945 140
rect 905 110 915 130
rect 935 110 945 130
rect 905 100 945 110
rect 725 90 945 100
rect 725 70 735 90
rect 755 70 915 90
rect 935 70 945 90
rect 725 60 945 70
rect 725 50 765 60
rect 725 30 735 50
rect 755 30 765 50
rect 725 20 765 30
rect 905 50 945 60
rect 905 30 915 50
rect 935 30 945 50
rect 905 20 945 30
rect 1205 -75 1245 145
rect 1275 85 1315 95
rect 1275 65 1285 85
rect 1305 65 1315 85
rect 1275 45 1315 65
rect 1275 25 1285 45
rect 1305 25 1315 45
rect 1275 -75 1315 25
rect -270 -385 -230 -370
rect -270 -405 -260 -385
rect -240 -405 -230 -385
rect -270 -420 -230 -405
rect 760 -400 900 -385
rect 760 -420 795 -400
rect 815 -420 840 -400
rect 860 -420 900 -400
rect 760 -435 900 -420
rect 1115 -400 1155 -385
rect 1115 -420 1125 -400
rect 1145 -420 1155 -400
rect 1115 -435 1155 -420
rect 210 -485 250 -470
rect 210 -505 220 -485
rect 240 -505 250 -485
rect 210 -520 250 -505
rect 650 -485 690 -470
rect 650 -505 660 -485
rect 680 -505 690 -485
rect 650 -520 690 -505
rect 320 -730 460 -715
rect 320 -750 355 -730
rect 375 -750 405 -730
rect 425 -750 460 -730
rect 320 -765 460 -750
rect -160 -830 95 -815
rect 370 -830 410 -765
rect -160 -850 -155 -830
rect -135 -850 -45 -830
rect -25 -850 95 -830
rect -160 -865 95 -850
rect 1225 -835 1365 -820
rect 1225 -855 1230 -835
rect 1250 -855 1340 -835
rect 1360 -855 1365 -835
rect 1225 -870 1365 -855
<< labels >>
rlabel metal1 -250 130 -250 130 5 B_M1
rlabel locali -180 0 -180 0 5 S_M1
rlabel locali -90 180 -90 180 1 D_M1
rlabel poly -135 -40 -135 -40 5 G_M1
rlabel metal1 125 135 125 135 5 B_M3
rlabel locali 195 0 195 0 1 S1_M3
rlabel locali 285 0 285 0 1 D1_M3
rlabel locali 375 0 375 0 1 S2_M3
rlabel locali 465 0 465 0 1 D2_M3
rlabel poly 330 -40 330 -40 1 G_M3
rlabel metal1 655 160 655 160 7 B_M4
rlabel locali 745 180 745 180 1 S1_M4
rlabel locali 835 180 835 180 1 D1_M4
rlabel locali 925 180 925 180 1 S2_M4
rlabel locali 1015 180 1015 180 1 D2_M4
rlabel metal1 880 270 880 270 1 G_M4
rlabel metal1 1225 180 1225 180 1 B_M2
rlabel locali 1295 175 1295 175 1 S_M2
rlabel locali 1385 175 1385 175 1 D_M2
rlabel poly 1340 -45 1340 -45 5 G_M2
rlabel metal1 -250 -420 -250 -420 5 B_M7
rlabel locali -180 -775 -180 -775 5 S1_M7
rlabel locali -90 -775 -90 -775 5 D_M7
rlabel locali 0 -775 0 -775 5 S2_M7
rlabel metal1 -90 -865 -90 -865 5 G_M7
rlabel locali 300 -475 300 -475 1 S_M8
rlabel locali 390 -675 390 -675 5 D_M8
rlabel locali 480 -475 480 -475 1 S2_M8
rlabel metal1 355 -765 355 -765 5 G_M8
rlabel metal1 1135 -435 1135 -435 5 B_M5
rlabel locali 1295 -380 1295 -380 1 D_M5
rlabel locali 1385 -780 1385 -780 5 S2_M5
rlabel metal1 1255 -870 1255 -870 5 G_M5
rlabel metal1 210 -485 210 -485 7 B_M8
rlabel locali 1205 -780 1205 -780 5 S1_M5
rlabel metal1 670 -485 670 -485 1 B_M6
rlabel locali 740 -675 740 -675 5 S1_M6
rlabel locali 830 -475 830 -475 1 D_M6
rlabel locali 920 -675 920 -675 5 S2_M6
rlabel metal1 825 -385 825 -385 1 G_M6
<< end >>
