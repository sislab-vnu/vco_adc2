magic
tech sky130A
timestamp 1726044335
<< nwell >>
rect -130 -40 300 340
<< pwell >>
rect -130 -350 300 -70
<< nmos >>
rect 0 -310 100 -110
rect 140 -310 240 -110
<< pmos >>
rect 0 0 100 300
rect 140 0 240 300
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -310 0 -300
rect 100 -120 140 -110
rect 100 -140 110 -120
rect 130 -140 140 -120
rect 100 -160 140 -140
rect 100 -180 110 -160
rect 130 -180 140 -160
rect 100 -200 140 -180
rect 100 -220 110 -200
rect 130 -220 140 -200
rect 100 -240 140 -220
rect 100 -260 110 -240
rect 130 -260 140 -240
rect 100 -280 140 -260
rect 100 -300 110 -280
rect 130 -300 140 -280
rect 100 -310 140 -300
rect 240 -120 280 -110
rect 240 -140 250 -120
rect 270 -140 280 -120
rect 240 -160 280 -140
rect 240 -180 250 -160
rect 270 -180 280 -160
rect 240 -200 280 -180
rect 240 -220 250 -200
rect 270 -220 280 -200
rect 240 -240 280 -220
rect 240 -260 250 -240
rect 270 -260 280 -240
rect 240 -280 280 -260
rect 240 -300 250 -280
rect 270 -300 280 -280
rect 240 -310 280 -300
<< pdiff >>
rect -40 290 0 300
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 100 290 140 300
rect 100 270 110 290
rect 130 270 140 290
rect 100 250 140 270
rect 100 230 110 250
rect 130 230 140 250
rect 100 210 140 230
rect 100 190 110 210
rect 130 190 140 210
rect 100 170 140 190
rect 100 150 110 170
rect 130 150 140 170
rect 100 130 140 150
rect 100 110 110 130
rect 130 110 140 130
rect 100 90 140 110
rect 100 70 110 90
rect 130 70 140 90
rect 100 50 140 70
rect 100 30 110 50
rect 130 30 140 50
rect 100 0 140 30
rect 240 290 280 300
rect 240 270 250 290
rect 270 270 280 290
rect 240 250 280 270
rect 240 230 250 250
rect 270 230 280 250
rect 240 210 280 230
rect 240 190 250 210
rect 270 190 280 210
rect 240 170 280 190
rect 240 150 250 170
rect 270 150 280 170
rect 240 130 280 150
rect 240 110 250 130
rect 270 110 280 130
rect 240 90 280 110
rect 240 70 250 90
rect 270 70 280 90
rect 240 50 280 70
rect 240 30 250 50
rect 270 30 280 50
rect 240 0 280 30
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect 110 -140 130 -120
rect 110 -180 130 -160
rect 110 -220 130 -200
rect 110 -260 130 -240
rect 110 -300 130 -280
rect 250 -140 270 -120
rect 250 -180 270 -160
rect 250 -220 270 -200
rect 250 -260 270 -240
rect 250 -300 270 -280
<< pdiffc >>
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 110 270 130 290
rect 110 230 130 250
rect 110 190 130 210
rect 110 150 130 170
rect 110 110 130 130
rect 110 70 130 90
rect 110 30 130 50
rect 250 270 270 290
rect 250 230 270 250
rect 250 190 270 210
rect 250 150 270 170
rect 250 110 270 130
rect 250 70 270 90
rect 250 30 270 50
<< psubdiff >>
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< nsubdiff >>
rect -110 290 -70 305
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
<< psubdiffcont >>
rect -100 -300 -80 -280
<< nsubdiffcont >>
rect -100 270 -80 290
<< poly >>
rect 0 300 100 340
rect 140 300 240 340
rect 0 -40 100 0
rect 140 -40 240 0
rect 0 -45 240 -40
rect 0 -65 35 -45
rect 55 -65 180 -45
rect 200 -65 240 -45
rect 0 -70 240 -65
rect 0 -110 100 -70
rect 140 -110 240 -70
rect 0 -350 100 -310
rect 140 -350 240 -310
<< polycont >>
rect 35 -65 55 -45
rect 180 -65 200 -45
<< locali >>
rect -40 390 280 430
rect -110 290 -70 305
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
rect -40 290 0 390
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 100 290 140 300
rect 100 270 110 290
rect 130 270 140 290
rect 100 250 140 270
rect 100 230 110 250
rect 130 230 140 250
rect 100 210 140 230
rect 100 190 110 210
rect 130 190 140 210
rect 100 170 140 190
rect 100 150 110 170
rect 130 150 140 170
rect 100 130 140 150
rect 100 110 110 130
rect 130 110 140 130
rect 100 90 140 110
rect 100 70 110 90
rect 130 70 140 90
rect 100 50 140 70
rect 100 30 110 50
rect 130 30 140 50
rect 25 -45 70 -35
rect 25 -65 35 -45
rect 55 -65 70 -45
rect 25 -80 70 -65
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -400 0 -300
rect 100 -120 140 30
rect 240 290 280 390
rect 240 270 250 290
rect 270 270 280 290
rect 240 250 280 270
rect 240 230 250 250
rect 270 230 280 250
rect 240 210 280 230
rect 240 190 250 210
rect 270 190 280 210
rect 240 170 280 190
rect 240 150 250 170
rect 270 150 280 170
rect 240 130 280 150
rect 240 110 250 130
rect 270 110 280 130
rect 240 90 280 110
rect 240 70 250 90
rect 270 70 280 90
rect 240 50 280 70
rect 240 30 250 50
rect 270 30 280 50
rect 240 0 280 30
rect 165 -45 210 -35
rect 165 -65 180 -45
rect 200 -65 210 -45
rect 165 -80 210 -65
rect 100 -140 110 -120
rect 130 -140 140 -120
rect 100 -160 140 -140
rect 100 -180 110 -160
rect 130 -180 140 -160
rect 100 -200 140 -180
rect 100 -220 110 -200
rect 130 -220 140 -200
rect 100 -240 140 -220
rect 100 -260 110 -240
rect 130 -260 140 -240
rect 100 -280 140 -260
rect 100 -300 110 -280
rect 130 -300 140 -280
rect 100 -310 140 -300
rect 240 -120 280 -110
rect 240 -140 250 -120
rect 270 -140 280 -120
rect 240 -160 280 -140
rect 240 -180 250 -160
rect 270 -180 280 -160
rect 240 -200 280 -180
rect 240 -220 250 -200
rect 270 -220 280 -200
rect 240 -240 280 -220
rect 240 -260 250 -240
rect 270 -260 280 -240
rect 240 -280 280 -260
rect 240 -300 250 -280
rect 270 -300 280 -280
rect 240 -400 280 -300
rect -40 -440 280 -400
<< viali >>
rect -100 270 -80 290
rect 35 -65 55 -45
rect -100 -300 -80 -280
rect 180 -65 200 -45
<< metal1 >>
rect -110 290 -70 305
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
rect 25 -45 210 -35
rect 25 -65 35 -45
rect 55 -65 180 -45
rect 200 -65 210 -45
rect 25 -80 210 -65
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< labels >>
rlabel locali 120 430 120 430 1 VPWR
port 1 n
rlabel metal1 -90 305 -90 305 1 VCCA
port 2 n
rlabel locali 120 300 120 300 1 Y
port 3 n
rlabel metal1 -90 -265 -90 -265 1 GND
port 4 n
rlabel locali 120 -400 120 -400 1 VGND
port 5 n
rlabel metal1 25 -55 25 -55 7 A
port 6 w
<< end >>
