magic
tech sky130A
magscale 1 2
timestamp 1729593089
<< nwell >>
rect 5530 2900 5770 3220
<< pwell >>
rect 5614 2684 5746 2836
<< psubdiff >>
rect 5640 2777 5720 2810
rect 5640 2743 5663 2777
rect 5697 2743 5720 2777
rect 5640 2710 5720 2743
<< nsubdiff >>
rect 5640 3077 5720 3110
rect 5640 3043 5663 3077
rect 5697 3043 5720 3077
rect 5640 3010 5720 3043
<< psubdiffcont >>
rect 5663 2743 5697 2777
<< nsubdiffcont >>
rect 5663 3043 5697 3077
<< locali >>
rect 780 6950 1660 7030
rect 19410 7010 19930 7030
rect 19410 6970 19440 7010
rect 19480 6970 19930 7010
rect 19410 6950 19930 6970
rect 5390 3890 5470 3900
rect 5390 3810 6850 3890
rect 5390 3800 5470 3810
rect 6850 3480 7040 3600
rect 5640 3077 5720 3110
rect 5640 3043 5663 3077
rect 5697 3043 5720 3077
rect 5640 3010 5720 3043
rect 4990 2910 5150 2970
rect 5560 2950 5610 2970
rect 5540 2947 5610 2950
rect 5540 2913 5543 2947
rect 5577 2913 5610 2947
rect 5540 2910 5610 2913
rect 5560 2870 5610 2910
rect 5640 2777 5720 2810
rect 5640 2743 5663 2777
rect 5697 2743 5720 2777
rect 5640 2710 5720 2743
<< viali >>
rect 5663 3043 5697 3077
rect 5543 2913 5577 2947
rect 5510 2740 5544 2774
rect 5663 2743 5697 2777
<< metal1 >>
rect 640 7230 1160 7330
rect 19310 7230 19930 7330
rect 4090 3790 4170 3900
rect 5110 3370 5950 3470
rect 5130 3230 5230 3370
rect 5640 3077 5720 3370
rect 5640 3043 5663 3077
rect 5697 3043 5720 3077
rect 5640 3010 5720 3043
rect 5490 2947 5610 2990
rect 5490 2913 5543 2947
rect 5577 2930 5610 2947
rect 5850 2930 5950 3370
rect 5577 2913 5950 2930
rect 5490 2870 5950 2913
rect 5480 2800 5570 2820
rect 4890 2774 5570 2800
rect 4890 2740 5510 2774
rect 5544 2740 5570 2774
rect 4890 2230 4990 2740
rect 5480 2730 5570 2740
rect 5640 2780 5720 2810
rect 6230 2780 6330 4200
rect 8230 3480 8410 3590
rect 5640 2777 6330 2780
rect 5640 2743 5663 2777
rect 5697 2743 6330 2777
rect 5640 2720 6330 2743
rect 5640 2710 5720 2720
rect 6230 2650 6330 2720
rect 5570 2590 6330 2650
rect 6310 2150 6600 2200
rect 5940 880 6640 980
rect 8400 0 8700 100
use sky130_fd_pr__res_generic_po_DKCPUZ  sky130_fd_pr__res_generic_po_DKCPUZ_0
timestamp 1729593089
transform 0 -1 4780 1 0 3848
box -48 -630 48 630
use sky130_fd_pr__res_generic_po_DKCPUZ  sky130_fd_pr__res_generic_po_DKCPUZ_1
timestamp 1729593089
transform 0 -1 7640 1 0 3538
box -48 -630 48 630
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0
timestamp 1729593089
transform 1 0 5128 0 1 2638
box -38 -48 498 592
use vco_ring_osc  vco_ring_osc_0
timestamp 1729593089
transform 1 0 600 0 1 4200
box -600 -4200 20040 3130
<< labels >>
rlabel metal1 s 5160 3470 5160 3470 4 VCCD
rlabel locali s 5020 2970 5020 2970 4 ENB
rlabel metal1 s 6470 980 6470 980 4 p[4]
rlabel metal1 s 4100 3900 4100 3900 4 Anlg_in
rlabel metal1 s 19900 7330 19900 7330 4 VCCA
rlabel locali s 19900 7030 19900 7030 4 VPWR
rlabel metal1 s 6230 3340 6230 3340 4 GND
<< end >>
