magic
tech sky130A
timestamp 1726544869
<< nwell >>
rect -130 -40 290 220
<< pmoshvt >>
rect 0 0 50 180
rect 90 0 140 180
rect 180 0 230 180
<< pdiff >>
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 70 0 110
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 70 90 110
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 170 180 180
rect 140 150 150 170
rect 170 150 180 170
rect 140 130 180 150
rect 140 110 150 130
rect 170 110 180 130
rect 140 70 180 110
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
rect 230 170 270 180
rect 230 150 240 170
rect 260 150 270 170
rect 230 130 270 150
rect 230 110 240 130
rect 260 110 270 130
rect 230 70 270 110
rect 230 50 240 70
rect 260 50 270 70
rect 230 30 270 50
rect 230 10 240 30
rect 260 10 270 30
rect 230 0 270 10
<< pdiffc >>
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 50 -10 70
rect -30 10 -10 30
rect 60 150 80 170
rect 60 110 80 130
rect 60 50 80 70
rect 60 10 80 30
rect 150 150 170 170
rect 150 110 170 130
rect 150 50 170 70
rect 150 10 170 30
rect 240 150 260 170
rect 240 110 260 130
rect 240 50 260 70
rect 240 10 260 30
<< nsubdiff >>
rect -110 170 -70 185
rect -110 150 -100 170
rect -80 150 -70 170
rect -110 135 -70 150
<< nsubdiffcont >>
rect -100 150 -80 170
<< poly >>
rect 0 250 230 260
rect 0 230 45 250
rect 65 230 105 250
rect 125 230 165 250
rect 185 230 230 250
rect 0 220 230 230
rect 0 180 50 220
rect 90 180 140 220
rect 180 180 230 220
rect 0 -40 50 0
rect 90 -40 140 0
rect 180 -40 230 0
<< polycont >>
rect 45 230 65 250
rect 105 230 125 250
rect 165 230 185 250
<< locali >>
rect 25 250 205 260
rect 25 230 45 250
rect 65 230 105 250
rect 125 230 165 250
rect 185 230 205 250
rect 25 220 205 230
rect -110 170 -70 185
rect -110 150 -100 170
rect -80 150 -70 170
rect -110 135 -70 150
rect -40 170 0 180
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 70 0 110
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 170 90 180
rect 50 150 60 170
rect 80 150 90 170
rect 50 130 90 150
rect 50 110 60 130
rect 80 110 90 130
rect 50 70 90 110
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 170 180 180
rect 140 150 150 170
rect 170 150 180 170
rect 140 130 180 150
rect 140 110 150 130
rect 170 110 180 130
rect 140 70 180 110
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
rect 230 170 270 180
rect 230 150 240 170
rect 260 150 270 170
rect 230 130 270 150
rect 230 110 240 130
rect 260 110 270 130
rect 230 70 270 110
rect 230 50 240 70
rect 260 50 270 70
rect 230 30 270 50
rect 230 10 240 30
rect 260 10 270 30
rect 230 0 270 10
<< viali >>
rect 45 230 65 250
rect 105 230 125 250
rect 165 230 185 250
rect -100 150 -80 170
rect -30 150 -10 170
rect -30 110 -10 130
rect 60 50 80 70
rect 60 10 80 30
rect 150 150 170 170
rect 150 110 170 130
rect 240 50 260 70
rect 240 10 260 30
<< metal1 >>
rect 0 250 230 260
rect 0 230 45 250
rect 65 230 105 250
rect 125 230 165 250
rect 185 230 230 250
rect 0 220 230 230
rect -110 170 -70 185
rect -110 150 -100 170
rect -80 150 -70 170
rect -110 135 -70 150
rect -40 170 0 180
rect -40 150 -30 170
rect -10 165 0 170
rect 140 170 180 180
rect 140 165 150 170
rect -10 150 150 165
rect 170 150 180 170
rect -40 130 180 150
rect -40 110 -30 130
rect -10 115 150 130
rect -10 110 0 115
rect -40 100 0 110
rect 140 110 150 115
rect 170 110 180 130
rect 140 100 180 110
rect 50 70 90 80
rect 50 50 60 70
rect 80 65 90 70
rect 230 70 270 80
rect 230 65 240 70
rect 80 50 240 65
rect 260 50 270 70
rect 50 30 270 50
rect 50 10 60 30
rect 80 15 240 30
rect 80 10 90 15
rect 50 0 90 10
rect 230 10 240 15
rect 260 10 270 30
rect 230 0 270 10
<< labels >>
rlabel metal1 -90 185 -90 185 1 B
rlabel metal1 -20 180 -20 180 1 S
rlabel metal1 250 0 250 0 5 D
rlabel metal1 115 260 115 260 5 G
<< end >>
