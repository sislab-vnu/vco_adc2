magic
tech sky130A
timestamp 1726718672
<< dnwell >>
rect 120 -1090 760 -460
rect 1970 -1110 2610 -480
<< nwell >>
rect 1555 215 1595 225
rect 1015 90 1035 110
rect 75 -565 805 -415
rect -1330 -860 -1170 -630
rect -1325 -885 -1170 -860
rect -1330 -910 -1170 -885
rect 75 -985 225 -565
rect 655 -985 805 -565
rect 75 -1140 805 -985
rect 1925 -585 2655 -435
rect 1925 -1005 2075 -585
rect 2505 -1005 2655 -585
rect 1925 -1155 2655 -1005
<< pwell >>
rect -1450 -870 -1360 -625
<< pdiffc >>
rect 1015 90 1035 110
<< psubdiff >>
rect -1430 -800 -1380 -790
rect -1430 -820 -1415 -800
rect -1395 -820 -1380 -800
rect -1430 -830 -1380 -820
<< nsubdiff >>
rect 95 -445 785 -435
rect 95 -465 135 -445
rect 155 -465 195 -445
rect 215 -465 255 -445
rect 275 -465 315 -445
rect 335 -465 375 -445
rect 395 -465 435 -445
rect 455 -465 495 -445
rect 515 -465 555 -445
rect 575 -465 615 -445
rect 635 -465 675 -445
rect 695 -465 735 -445
rect 755 -465 785 -445
rect 95 -475 785 -465
rect 95 -515 135 -475
rect 95 -535 110 -515
rect 130 -535 135 -515
rect 95 -575 135 -535
rect 95 -595 110 -575
rect 130 -595 135 -575
rect 95 -635 135 -595
rect 95 -655 110 -635
rect 130 -655 135 -635
rect 95 -695 135 -655
rect 95 -715 110 -695
rect 130 -715 135 -695
rect 95 -755 135 -715
rect 95 -775 110 -755
rect 130 -775 135 -755
rect -1270 -800 -1220 -790
rect -1270 -820 -1255 -800
rect -1235 -820 -1220 -800
rect -1270 -830 -1220 -820
rect 95 -815 135 -775
rect 95 -835 110 -815
rect 130 -835 135 -815
rect 95 -875 135 -835
rect 95 -895 110 -875
rect 130 -895 135 -875
rect 95 -935 135 -895
rect 95 -955 110 -935
rect 130 -955 135 -935
rect 95 -995 135 -955
rect 95 -1015 110 -995
rect 130 -1015 135 -995
rect 95 -1055 135 -1015
rect 95 -1075 110 -1055
rect 130 -1075 135 -1055
rect 745 -485 785 -475
rect 745 -505 755 -485
rect 775 -505 785 -485
rect 745 -545 785 -505
rect 745 -565 755 -545
rect 775 -565 785 -545
rect 745 -605 785 -565
rect 745 -625 755 -605
rect 775 -625 785 -605
rect 745 -665 785 -625
rect 745 -685 755 -665
rect 775 -685 785 -665
rect 745 -725 785 -685
rect 745 -745 755 -725
rect 775 -745 785 -725
rect 745 -785 785 -745
rect 745 -805 755 -785
rect 775 -805 785 -785
rect 745 -845 785 -805
rect 745 -865 755 -845
rect 775 -865 785 -845
rect 745 -905 785 -865
rect 745 -925 755 -905
rect 775 -925 785 -905
rect 745 -965 785 -925
rect 745 -985 755 -965
rect 775 -985 785 -965
rect 745 -1025 785 -985
rect 745 -1045 755 -1025
rect 775 -1045 785 -1025
rect 745 -1075 785 -1045
rect 95 -1085 785 -1075
rect 95 -1105 150 -1085
rect 170 -1105 210 -1085
rect 230 -1105 270 -1085
rect 290 -1105 330 -1085
rect 350 -1105 390 -1085
rect 410 -1105 455 -1085
rect 475 -1105 515 -1085
rect 535 -1105 575 -1085
rect 595 -1105 635 -1085
rect 655 -1105 695 -1085
rect 715 -1105 755 -1085
rect 775 -1105 785 -1085
rect 95 -1120 785 -1105
rect 1945 -465 2635 -455
rect 1945 -485 1985 -465
rect 2005 -485 2045 -465
rect 2065 -485 2105 -465
rect 2125 -485 2165 -465
rect 2185 -485 2225 -465
rect 2245 -485 2285 -465
rect 2305 -485 2345 -465
rect 2365 -485 2405 -465
rect 2425 -485 2465 -465
rect 2485 -485 2525 -465
rect 2545 -485 2585 -465
rect 2605 -485 2635 -465
rect 1945 -495 2635 -485
rect 1945 -535 1985 -495
rect 1945 -555 1955 -535
rect 1975 -555 1985 -535
rect 1945 -595 1985 -555
rect 1945 -615 1955 -595
rect 1975 -615 1985 -595
rect 1945 -655 1985 -615
rect 1945 -675 1955 -655
rect 1975 -675 1985 -655
rect 1945 -715 1985 -675
rect 1945 -735 1955 -715
rect 1975 -735 1985 -715
rect 1945 -775 1985 -735
rect 1945 -795 1955 -775
rect 1975 -795 1985 -775
rect 1945 -835 1985 -795
rect 1945 -855 1955 -835
rect 1975 -855 1985 -835
rect 1945 -895 1985 -855
rect 1945 -915 1955 -895
rect 1975 -915 1985 -895
rect 1945 -955 1985 -915
rect 1945 -975 1955 -955
rect 1975 -975 1985 -955
rect 1945 -1015 1985 -975
rect 1945 -1035 1955 -1015
rect 1975 -1035 1985 -1015
rect 1945 -1075 1985 -1035
rect 1945 -1095 1955 -1075
rect 1975 -1095 1985 -1075
rect 2595 -505 2635 -495
rect 2595 -525 2605 -505
rect 2625 -525 2635 -505
rect 2595 -565 2635 -525
rect 2595 -585 2605 -565
rect 2625 -585 2635 -565
rect 2595 -625 2635 -585
rect 2595 -645 2605 -625
rect 2625 -645 2635 -625
rect 2595 -685 2635 -645
rect 2595 -705 2605 -685
rect 2625 -705 2635 -685
rect 2595 -745 2635 -705
rect 2595 -765 2605 -745
rect 2625 -765 2635 -745
rect 2595 -805 2635 -765
rect 2595 -825 2605 -805
rect 2625 -825 2635 -805
rect 2595 -865 2635 -825
rect 2595 -885 2605 -865
rect 2625 -885 2635 -865
rect 2595 -925 2635 -885
rect 2595 -945 2605 -925
rect 2625 -945 2635 -925
rect 2595 -985 2635 -945
rect 2595 -1005 2605 -985
rect 2625 -1005 2635 -985
rect 2595 -1045 2635 -1005
rect 2595 -1065 2605 -1045
rect 2625 -1065 2635 -1045
rect 2595 -1095 2635 -1065
rect 1945 -1100 2635 -1095
rect 1945 -1105 2605 -1100
rect 1945 -1125 1990 -1105
rect 2010 -1125 2050 -1105
rect 2070 -1125 2110 -1105
rect 2130 -1125 2170 -1105
rect 2190 -1125 2230 -1105
rect 2250 -1125 2290 -1105
rect 2310 -1125 2350 -1105
rect 2370 -1125 2410 -1105
rect 2430 -1125 2470 -1105
rect 2490 -1125 2530 -1105
rect 2550 -1120 2605 -1105
rect 2625 -1120 2635 -1100
rect 2550 -1125 2635 -1120
rect 1945 -1135 2635 -1125
<< psubdiffcont >>
rect -1415 -820 -1395 -800
<< nsubdiffcont >>
rect 135 -465 155 -445
rect 195 -465 215 -445
rect 255 -465 275 -445
rect 315 -465 335 -445
rect 375 -465 395 -445
rect 435 -465 455 -445
rect 495 -465 515 -445
rect 555 -465 575 -445
rect 615 -465 635 -445
rect 675 -465 695 -445
rect 735 -465 755 -445
rect 110 -535 130 -515
rect 110 -595 130 -575
rect 110 -655 130 -635
rect 110 -715 130 -695
rect 110 -775 130 -755
rect -1255 -820 -1235 -800
rect 110 -835 130 -815
rect 110 -895 130 -875
rect 110 -955 130 -935
rect 110 -1015 130 -995
rect 110 -1075 130 -1055
rect 755 -505 775 -485
rect 755 -565 775 -545
rect 755 -625 775 -605
rect 755 -685 775 -665
rect 755 -745 775 -725
rect 755 -805 775 -785
rect 755 -865 775 -845
rect 755 -925 775 -905
rect 755 -985 775 -965
rect 755 -1045 775 -1025
rect 150 -1105 170 -1085
rect 210 -1105 230 -1085
rect 270 -1105 290 -1085
rect 330 -1105 350 -1085
rect 390 -1105 410 -1085
rect 455 -1105 475 -1085
rect 515 -1105 535 -1085
rect 575 -1105 595 -1085
rect 635 -1105 655 -1085
rect 695 -1105 715 -1085
rect 755 -1105 775 -1085
rect 1985 -485 2005 -465
rect 2045 -485 2065 -465
rect 2105 -485 2125 -465
rect 2165 -485 2185 -465
rect 2225 -485 2245 -465
rect 2285 -485 2305 -465
rect 2345 -485 2365 -465
rect 2405 -485 2425 -465
rect 2465 -485 2485 -465
rect 2525 -485 2545 -465
rect 2585 -485 2605 -465
rect 1955 -555 1975 -535
rect 1955 -615 1975 -595
rect 1955 -675 1975 -655
rect 1955 -735 1975 -715
rect 1955 -795 1975 -775
rect 1955 -855 1975 -835
rect 1955 -915 1975 -895
rect 1955 -975 1975 -955
rect 1955 -1035 1975 -1015
rect 1955 -1095 1975 -1075
rect 2605 -525 2625 -505
rect 2605 -585 2625 -565
rect 2605 -645 2625 -625
rect 2605 -705 2625 -685
rect 2605 -765 2625 -745
rect 2605 -825 2625 -805
rect 2605 -885 2625 -865
rect 2605 -945 2625 -925
rect 2605 -1005 2625 -985
rect 2605 -1065 2625 -1045
rect 1990 -1125 2010 -1105
rect 2050 -1125 2070 -1105
rect 2110 -1125 2130 -1105
rect 2170 -1125 2190 -1105
rect 2230 -1125 2250 -1105
rect 2290 -1125 2310 -1105
rect 2350 -1125 2370 -1105
rect 2410 -1125 2430 -1105
rect 2470 -1125 2490 -1105
rect 2530 -1125 2550 -1105
rect 2605 -1120 2625 -1100
<< poly >>
rect 130 -10 180 0
rect 130 -30 145 -10
rect 165 -30 180 -10
rect 130 -40 180 -30
rect 1595 -10 1645 0
rect 1595 -30 1610 -10
rect 1630 -30 1645 -10
rect 1595 -40 1645 -30
<< polycont >>
rect 145 -30 165 -10
rect 1610 -30 1630 -10
<< locali >>
rect 90 415 495 455
rect 90 225 130 415
rect 455 225 495 415
rect 60 210 130 225
rect 60 175 90 210
rect 425 200 495 225
rect 425 175 455 200
rect 975 175 1005 220
rect 1525 215 1595 225
rect 1525 175 1555 215
rect 1645 100 1835 175
rect 130 -10 180 0
rect 130 -30 145 -10
rect 165 -30 180 -10
rect 130 -40 180 -30
rect 1095 -245 1135 40
rect 1595 -10 1645 0
rect 1595 -30 1610 -10
rect 1630 -30 1645 -10
rect 1595 -40 1645 -30
rect -1360 -470 -1325 -365
rect -895 -425 -185 -375
rect 3725 -400 3765 -250
rect -1355 -585 -1325 -570
rect -895 -580 -855 -425
rect -1350 -675 -1330 -585
rect -925 -595 -855 -580
rect -1355 -685 -1325 -675
rect -1355 -705 -1350 -685
rect -1330 -705 -1325 -685
rect -1430 -800 -1380 -790
rect -1430 -820 -1415 -800
rect -1395 -820 -1380 -800
rect -1430 -830 -1380 -820
rect -1355 -860 -1325 -705
rect -1220 -790 -1165 -625
rect -925 -630 -895 -595
rect -415 -705 -375 -425
rect 95 -445 785 -435
rect 95 -465 135 -445
rect 155 -465 195 -445
rect 215 -465 255 -445
rect 275 -465 315 -445
rect 335 -465 375 -445
rect 395 -465 435 -445
rect 455 -465 495 -445
rect 515 -465 555 -445
rect 575 -465 615 -445
rect 635 -465 675 -445
rect 695 -465 735 -445
rect 755 -465 785 -445
rect 3430 -450 4140 -400
rect 95 -475 785 -465
rect 95 -515 135 -475
rect 95 -535 110 -515
rect 130 -535 135 -515
rect 95 -575 135 -535
rect 95 -595 110 -575
rect 130 -595 135 -575
rect 95 -635 135 -595
rect 95 -655 110 -635
rect 130 -655 135 -635
rect 95 -695 135 -655
rect -1270 -800 -1165 -790
rect -1270 -820 -1255 -800
rect -1235 -820 -1205 -800
rect -1185 -820 -1165 -800
rect -1270 -830 -1165 -820
rect 95 -715 110 -695
rect 130 -715 135 -695
rect 95 -755 135 -715
rect 95 -775 110 -755
rect 130 -775 135 -755
rect 95 -815 135 -775
rect 95 -835 110 -815
rect 130 -835 135 -815
rect -1350 -885 -1330 -860
rect 95 -875 135 -835
rect 95 -895 110 -875
rect 130 -895 135 -875
rect -1355 -950 -1330 -945
rect -1350 -1010 -1330 -950
rect -1355 -1075 -1330 -1010
rect -1355 -1090 -1295 -1075
rect -1355 -1120 -1340 -1090
rect -1310 -1120 -1295 -1090
rect -1355 -1135 -1295 -1120
rect -805 -1160 -765 -980
rect -325 -1160 -285 -905
rect 95 -935 135 -895
rect 95 -955 110 -935
rect 130 -955 135 -935
rect 95 -995 135 -955
rect 95 -1015 110 -995
rect 130 -1015 135 -995
rect 95 -1055 135 -1015
rect 95 -1075 110 -1055
rect 130 -1075 135 -1055
rect 745 -485 785 -475
rect 745 -505 755 -485
rect 775 -505 785 -485
rect 745 -545 785 -505
rect 745 -565 755 -545
rect 775 -565 785 -545
rect 745 -605 785 -565
rect 745 -625 755 -605
rect 775 -625 785 -605
rect 745 -665 785 -625
rect 745 -685 755 -665
rect 775 -685 785 -665
rect 745 -725 785 -685
rect 745 -745 755 -725
rect 775 -745 785 -725
rect 745 -785 785 -745
rect 745 -805 755 -785
rect 775 -805 785 -785
rect 745 -845 785 -805
rect 745 -865 755 -845
rect 775 -865 785 -845
rect 745 -905 785 -865
rect 745 -925 755 -905
rect 775 -925 785 -905
rect 745 -965 785 -925
rect 745 -985 755 -965
rect 775 -985 785 -965
rect 745 -1025 785 -985
rect 745 -1045 755 -1025
rect 775 -1045 785 -1025
rect 745 -1075 785 -1045
rect 95 -1085 785 -1075
rect 95 -1105 150 -1085
rect 170 -1105 210 -1085
rect 230 -1105 270 -1085
rect 290 -1105 330 -1085
rect 350 -1105 390 -1085
rect 410 -1105 455 -1085
rect 475 -1105 515 -1085
rect 535 -1105 575 -1085
rect 595 -1105 635 -1085
rect 655 -1105 695 -1085
rect 715 -1105 755 -1085
rect 775 -1105 785 -1085
rect 95 -1120 785 -1105
rect 1945 -465 2635 -455
rect 1945 -485 1985 -465
rect 2005 -485 2045 -465
rect 2065 -485 2105 -465
rect 2125 -485 2165 -465
rect 2185 -485 2225 -465
rect 2245 -485 2285 -465
rect 2305 -485 2345 -465
rect 2365 -485 2405 -465
rect 2425 -485 2465 -465
rect 2485 -485 2525 -465
rect 2545 -485 2585 -465
rect 2605 -485 2635 -465
rect 1945 -495 2635 -485
rect 1945 -535 1985 -495
rect 1945 -555 1955 -535
rect 1975 -555 1985 -535
rect 1945 -595 1985 -555
rect 1945 -615 1955 -595
rect 1975 -615 1985 -595
rect 1945 -655 1985 -615
rect 1945 -675 1955 -655
rect 1975 -675 1985 -655
rect 1945 -715 1985 -675
rect 1945 -735 1955 -715
rect 1975 -735 1985 -715
rect 1945 -775 1985 -735
rect 1945 -795 1955 -775
rect 1975 -795 1985 -775
rect 1945 -835 1985 -795
rect 1945 -855 1955 -835
rect 1975 -855 1985 -835
rect 1945 -895 1985 -855
rect 1945 -915 1955 -895
rect 1975 -915 1985 -895
rect 1945 -955 1985 -915
rect 1945 -975 1955 -955
rect 1975 -975 1985 -955
rect 1945 -1015 1985 -975
rect 1945 -1035 1955 -1015
rect 1975 -1035 1985 -1015
rect 1945 -1075 1985 -1035
rect 1945 -1095 1955 -1075
rect 1975 -1095 1985 -1075
rect 2595 -505 2635 -495
rect 2595 -525 2605 -505
rect 2625 -525 2635 -505
rect 2595 -565 2635 -525
rect 2595 -585 2605 -565
rect 2625 -585 2635 -565
rect 2595 -625 2635 -585
rect 2595 -645 2605 -625
rect 2625 -645 2635 -625
rect 2595 -685 2635 -645
rect 2595 -705 2605 -685
rect 2625 -705 2635 -685
rect 2595 -745 2635 -705
rect 3660 -735 3700 -450
rect 4100 -605 4140 -450
rect 4070 -625 4140 -605
rect 4070 -655 4100 -625
rect 2595 -765 2605 -745
rect 2625 -765 2635 -745
rect 2595 -805 2635 -765
rect 2595 -825 2605 -805
rect 2625 -825 2635 -805
rect 2595 -865 2635 -825
rect 2595 -885 2605 -865
rect 2625 -885 2635 -865
rect 2595 -925 2635 -885
rect 2595 -945 2605 -925
rect 2625 -945 2635 -925
rect 2595 -985 2635 -945
rect 2595 -1005 2605 -985
rect 2625 -1005 2635 -985
rect 2595 -1045 2635 -1005
rect 2595 -1065 2605 -1045
rect 2625 -1065 2635 -1045
rect 2595 -1095 2635 -1065
rect 1945 -1100 2635 -1095
rect 1945 -1105 2605 -1100
rect 1945 -1125 1990 -1105
rect 2010 -1125 2050 -1105
rect 2070 -1125 2110 -1105
rect 2130 -1125 2170 -1105
rect 2190 -1125 2230 -1105
rect 2250 -1125 2290 -1105
rect 2310 -1125 2350 -1105
rect 2370 -1125 2410 -1105
rect 2430 -1125 2470 -1105
rect 2490 -1125 2530 -1105
rect 2550 -1120 2605 -1105
rect 2625 -1120 2635 -1100
rect 2550 -1125 2635 -1120
rect 1945 -1135 2635 -1125
rect -805 -1210 -285 -1160
rect 3750 -1185 3790 -930
rect 4190 -1185 4230 -1005
rect 4465 -1185 4515 -250
rect -805 -1240 -765 -1210
rect 3750 -1235 4515 -1185
rect 180 -1530 220 -1295
rect 180 -1565 295 -1530
rect 1345 -1565 1620 -1530
<< viali >>
rect 190 190 210 210
rect 1565 190 1585 210
rect 190 150 210 170
rect 1565 150 1585 170
rect 1015 90 1035 110
rect 1015 50 1035 70
rect 145 -30 165 -10
rect 1610 -30 1630 -10
rect -1350 -705 -1330 -685
rect -1415 -820 -1395 -800
rect -1255 -820 -1235 -800
rect -1205 -820 -1185 -800
rect -1340 -1120 -1310 -1090
<< metal1 >>
rect 180 335 1595 385
rect 180 210 220 335
rect 495 260 725 300
rect 1045 260 1275 300
rect 180 190 190 210
rect 210 190 220 210
rect 180 170 220 190
rect 180 150 190 170
rect 210 150 220 170
rect 180 140 220 150
rect 1555 210 1595 335
rect 1555 190 1565 210
rect 1585 190 1595 210
rect 1555 170 1595 190
rect 1555 150 1565 170
rect 1585 150 1595 170
rect 1555 140 1595 150
rect 1005 110 1045 120
rect 1005 105 1015 110
rect 765 90 1015 105
rect 1035 90 1045 110
rect 765 70 1045 90
rect 765 55 1015 70
rect 1005 50 1015 55
rect 1035 50 1045 70
rect 1005 40 1045 50
rect 130 -10 180 0
rect 130 -30 145 -10
rect 165 -30 180 -10
rect 130 -40 180 -30
rect 1595 -10 1645 0
rect 1595 -30 1610 -10
rect 1630 -30 1645 -10
rect 1595 -40 1645 -30
rect -1110 -320 -185 -270
rect -1485 -455 -1435 -420
rect -1485 -790 -1435 -635
rect -1360 -680 -1320 -675
rect -1110 -680 -1060 -320
rect -810 -510 -760 -320
rect 3430 -345 3510 -295
rect -1360 -685 -1060 -680
rect -1360 -705 -1350 -685
rect -1330 -705 -1060 -685
rect -1360 -710 -1060 -705
rect -1360 -715 -1320 -710
rect -1485 -800 -1380 -790
rect -1485 -820 -1415 -800
rect -1395 -820 -1380 -800
rect -1485 -830 -1380 -820
rect -1270 -800 -1165 -790
rect -1270 -820 -1255 -800
rect -1235 -820 -1205 -800
rect -1185 -820 -1165 -800
rect -1270 -830 -1165 -820
rect -1485 -870 -1435 -830
rect -1220 -870 -1165 -830
rect 3460 -970 3510 -345
rect 3915 -570 4140 -520
rect -415 -1075 -365 -985
rect 3460 -1010 3610 -970
rect -1355 -1090 -185 -1075
rect -1355 -1120 -1340 -1090
rect -1310 -1120 -185 -1090
rect 3915 -1100 3965 -570
rect -1355 -1135 -185 -1120
rect 3395 -1160 3965 -1100
use n_lk  n_lk_2
timestamp 1726647885
transform 1 0 405 0 1 -895
box -130 -40 200 280
use n_lk  n_lk_3
timestamp 1726647885
transform 1 0 2255 0 1 -915
box -130 -40 200 280
use p_br1  p_br1_0
timestamp 1726647752
transform 1 0 130 0 1 40
box -130 -40 108 220
use p_br1  p_br1_1
timestamp 1726647752
transform 1 0 1595 0 1 40
box -130 -40 108 220
use p_br2  p_br2_0
timestamp 1726647805
transform 1 0 495 0 1 40
box -130 -40 290 260
use p_br2  p_br2_1
timestamp 1726647805
transform 1 0 1045 0 1 40
box -130 -40 290 260
use p_lk  p_lk_0
timestamp 1726647848
transform 1 0 -855 0 1 -985
box -130 -40 200 490
use p_lk  p_lk_1
timestamp 1726647848
transform 1 0 4140 0 1 -1010
box -130 -40 200 490
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 ~/eda/unic-cass/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -1461 -1 0 -453
box -19 -24 203 296
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 ~/eda/unic-cass/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 0 1 -1461 -1 0 -868
box -19 -24 157 296
<< labels >>
rlabel metal1 220 385 220 385 1 note_12
rlabel metal1 850 105 850 105 1 note_34
rlabel locali 255 -1530 255 -1530 1 input_R
rlabel locali 130 455 130 455 1 VCCA
port 1 n
rlabel metal1 155 -40 155 -40 5 Vbs1
port 3 s
rlabel metal1 1620 -40 1620 -40 5 Vbs2
port 4 s
rlabel metal1 610 300 610 300 1 Vbs3
rlabel metal1 565 300 565 300 1 Vbs3
port 5 n
rlabel metal1 1100 300 1100 300 1 Vbs4
port 6 n
rlabel locali 3700 -400 3700 -400 1 add_pwr
rlabel locali -1340 -365 -1340 -365 1 Dctrl
port 2 n
rlabel metal1 -1130 -680 -1130 -680 1 Open
rlabel metal1 -1120 -1075 -1120 -1075 1 lock
rlabel metal1 -1485 -430 -1485 -430 7 gnd
<< end >>
