magic
tech sky130A
timestamp 1730442989
<< nwell >>
rect 375 985 395 1005
rect -45 925 130 975
rect 1645 905 1865 1025
rect 1900 925 1905 975
rect 2415 825 2435 845
rect 2415 785 2435 805
<< pwell >>
rect 2415 340 2435 360
rect 2415 300 2435 320
<< polycont >>
rect 1075 570 1095 590
rect 1115 570 1135 590
rect 1155 570 1175 590
rect 1560 570 1580 590
rect 1600 570 1620 590
rect 1640 570 1660 590
<< locali >>
rect 805 1225 2095 1265
rect 910 1135 950 1225
rect 1455 1135 1495 1225
rect 1065 605 1185 615
rect 1550 610 1670 615
rect 650 590 1185 605
rect 650 570 1075 590
rect 1095 570 1115 590
rect 1135 570 1155 590
rect 1175 570 1185 590
rect 650 555 1185 570
rect 1355 590 1670 610
rect 1355 570 1560 590
rect 1580 570 1600 590
rect 1620 570 1640 590
rect 1660 570 1670 590
rect 1355 560 1670 570
rect 650 495 700 555
rect 1065 550 1185 555
rect 1550 550 1670 560
rect 405 445 700 495
rect 910 40 950 130
rect 1455 40 1495 130
rect 810 0 2000 40
<< viali >>
rect 375 985 395 1005
rect 1870 985 1890 1005
rect 375 945 395 965
rect 1870 945 1890 965
rect 375 905 395 925
rect 1870 905 1890 925
rect 1325 825 1345 845
rect 2415 825 2435 845
rect 1325 785 1345 805
rect 2415 785 2435 805
rect 1325 745 1345 765
rect 2415 745 2435 765
rect 1075 570 1095 590
rect 1115 570 1135 590
rect 1155 570 1175 590
rect 1560 570 1580 590
rect 1600 570 1620 590
rect 1640 570 1660 590
rect 2415 340 2435 360
rect 2415 300 2435 320
rect 2415 260 2435 280
<< metal1 >>
rect -110 1365 1970 1415
rect -110 1140 -70 1365
rect 840 1140 880 1365
rect 1385 1140 1425 1365
rect 1930 1140 1970 1365
rect 365 1005 405 1025
rect 365 985 375 1005
rect 395 985 405 1005
rect 365 975 405 985
rect 1860 1005 1900 1025
rect 1860 985 1870 1005
rect 1890 985 1900 1005
rect 1860 975 1900 985
rect -130 925 270 975
rect 220 615 270 925
rect 365 965 2870 975
rect 365 945 375 965
rect 395 945 1870 965
rect 1890 945 2870 965
rect 365 925 2870 945
rect 365 905 375 925
rect 395 905 405 925
rect 365 885 405 905
rect 1100 615 1150 925
rect 1860 905 1870 925
rect 1890 905 1900 925
rect 1860 885 1900 905
rect 1315 845 1355 855
rect 1315 825 1325 845
rect 1345 825 1355 845
rect 1315 820 1355 825
rect 2405 845 2445 855
rect 2405 825 2415 845
rect 2435 825 2445 845
rect 2405 820 2445 825
rect 1315 805 2445 820
rect 1315 785 1325 805
rect 1345 785 2415 805
rect 2435 785 2445 805
rect 1315 770 2445 785
rect 1315 765 1355 770
rect 1315 745 1325 765
rect 1345 745 1355 765
rect 1315 735 1355 745
rect 1585 615 1635 770
rect 2405 765 2445 770
rect 2405 745 2415 765
rect 2435 745 2445 765
rect 2405 735 2445 745
rect 1065 590 1185 615
rect 1065 570 1075 590
rect 1095 570 1115 590
rect 1135 570 1155 590
rect 1175 570 1185 590
rect 1065 550 1185 570
rect 1550 590 1670 615
rect 1550 570 1560 590
rect 1580 570 1600 590
rect 1620 570 1640 590
rect 1660 570 1670 590
rect 1550 550 1670 570
rect 2035 555 2120 605
rect 2035 340 2085 555
rect -130 290 2085 340
rect 2405 360 2445 370
rect 2405 340 2415 360
rect 2435 340 2445 360
rect 2405 320 2870 340
rect 2405 300 2415 320
rect 2435 300 2870 320
rect 2405 290 2870 300
rect 2405 280 2445 290
rect 2405 260 2415 280
rect 2435 260 2445 280
rect 2405 250 2445 260
rect -110 -100 -70 125
rect 840 -100 880 125
rect 1385 -100 1425 125
rect 1930 -100 1970 125
rect -110 -150 1970 -100
use vco_aux_inv  vco_aux_inv_0
timestamp 1729846784
transform 1 0 950 0 1 640
box -130 -550 425 535
use vco_aux_inv  vco_aux_inv_1
timestamp 1729846784
transform 1 0 1495 0 1 640
box -130 -550 425 535
use vco_main_inv  vco_main_inv_0
timestamp 1730431575
transform 1 0 0 0 1 635
box -130 -635 830 630
use vco_main_inv  vco_main_inv_1
timestamp 1730431575
transform 1 0 2040 0 1 635
box -130 -635 830 630
<< labels >>
rlabel locali 1415 1265 1415 1265 1 VPWR
port 3 n
rlabel locali 1415 0 1415 0 5 VGND
port 4 s
rlabel metal1 -90 1415 -90 1415 1 VCCA
port 7 n
rlabel metal1 -95 -150 -95 -150 5 GND
port 8 s
rlabel metal1 -130 950 -130 950 7 inp
port 1 w
rlabel metal1 -130 310 -130 310 7 inn
port 2 w
rlabel metal1 2870 950 2870 950 3 outp
port 5 e
rlabel metal1 2870 310 2870 310 3 outn
port 6 e
<< end >>
