magic
tech sky130A
timestamp 1726913973
<< nwell >>
rect -145 -385 -25 -220
rect 975 -390 1125 -220
rect -185 -910 -100 -745
rect 805 -955 905 -790
rect -95 -1420 -10 -1410
rect 980 -1415 1175 -1410
rect -95 -1570 -20 -1420
rect 980 -1570 1140 -1415
rect -95 -1575 -10 -1570
rect 980 -1575 1175 -1570
<< pwell >>
rect -430 -505 -345 -435
rect -165 -505 -5 -435
rect 920 -505 1145 -435
rect -200 -1025 -100 -935
rect 785 -1075 925 -1005
rect -115 -1385 35 -1290
rect 960 -1360 1160 -1290
<< psubdiff >>
rect -410 -455 -370 -440
rect -410 -475 -400 -455
rect -380 -475 -370 -455
rect -410 -490 -370 -475
rect -165 -965 -125 -950
rect -165 -985 -155 -965
rect -135 -985 -125 -965
rect -165 -1000 -125 -985
rect 830 -1030 880 -1020
rect 830 -1050 845 -1030
rect 865 -1050 880 -1030
rect 830 -1060 880 -1050
rect 1020 -1315 1070 -1305
rect 1020 -1335 1035 -1315
rect 1055 -1335 1070 -1315
rect 1020 -1345 1070 -1335
<< nsubdiff >>
rect -105 -295 -65 -280
rect -105 -315 -95 -295
rect -75 -315 -65 -295
rect -105 -330 -65 -315
rect -165 -820 -125 -805
rect -165 -840 -155 -820
rect -135 -840 -125 -820
rect -165 -855 -125 -840
rect 840 -875 880 -860
rect 840 -895 850 -875
rect 870 -895 880 -875
rect 840 -910 880 -895
rect -65 -1470 -25 -1455
rect -65 -1490 -55 -1470
rect -35 -1490 -25 -1470
rect -65 -1505 -25 -1490
<< psubdiffcont >>
rect -400 -475 -380 -455
rect -155 -985 -135 -965
rect 845 -1050 865 -1030
rect 1035 -1335 1055 -1315
<< nsubdiffcont >>
rect -95 -315 -75 -295
rect -155 -840 -135 -820
rect 850 -895 870 -875
rect -55 -1490 -35 -1470
<< locali >>
rect -175 -255 -5 -220
rect -105 -295 -65 -255
rect 955 -270 1140 -220
rect -105 -315 -95 -295
rect -75 -315 -65 -295
rect -105 -330 -65 -315
rect -220 -405 10 -385
rect 910 -390 1150 -380
rect 910 -410 1050 -390
rect 1070 -410 1150 -390
rect 910 -420 1150 -410
rect -410 -455 -370 -440
rect -410 -475 -400 -455
rect -380 -475 -370 -455
rect -410 -490 -370 -475
rect -175 -491 -120 -490
rect -70 -491 -5 -490
rect -175 -540 -5 -491
rect 955 -540 1140 -495
rect -165 -820 -125 -805
rect -165 -840 -155 -820
rect -135 -840 -125 -820
rect -165 -855 -125 -840
rect 840 -875 880 -860
rect 840 -895 850 -875
rect 870 -895 880 -875
rect 840 -910 880 -895
rect 730 -950 900 -945
rect -165 -965 -125 -950
rect -165 -985 -155 -965
rect -135 -985 -125 -965
rect 730 -970 935 -950
rect -165 -1000 -125 -985
rect 830 -1030 880 -1020
rect 830 -1050 845 -1030
rect 865 -1050 880 -1030
rect 830 -1060 880 -1050
rect 1020 -1315 1070 -1305
rect 1020 -1335 1035 -1315
rect 1055 -1335 1070 -1315
rect 1020 -1345 1070 -1335
rect -124 -1413 53 -1389
rect -65 -1470 -25 -1455
rect -65 -1490 -55 -1470
rect -35 -1490 -25 -1470
rect -65 -1505 -25 -1490
<< viali >>
rect -95 -315 -75 -295
rect 180 -395 200 -375
rect 1050 -410 1070 -390
rect -400 -475 -380 -455
rect -155 -840 -135 -820
rect 850 -895 870 -875
rect -319 -927 -299 -907
rect -155 -985 -135 -965
rect 512 -976 529 -959
rect 569 -975 586 -958
rect 845 -1050 865 -1030
rect 1035 -1335 1055 -1315
rect 46 -1357 66 -1337
rect -55 -1490 -35 -1470
<< metal1 >>
rect -105 -295 -65 -280
rect -105 -315 -95 -295
rect -75 -315 -65 -295
rect -105 -330 -65 -315
rect -105 -375 210 -365
rect -105 -395 180 -375
rect 200 -395 210 -375
rect -105 -405 210 -395
rect 1040 -390 1075 -380
rect -410 -455 -370 -440
rect -410 -475 -400 -455
rect -380 -475 -370 -455
rect -410 -490 -370 -475
rect -105 -570 -70 -405
rect 1040 -410 1050 -390
rect 1070 -410 1075 -390
rect 1040 -665 1075 -410
rect 305 -700 1075 -665
rect -165 -820 -125 -805
rect -165 -840 -155 -820
rect -135 -840 -125 -820
rect -165 -855 -125 -840
rect 305 -865 340 -700
rect 305 -900 595 -865
rect -415 -907 -290 -900
rect -415 -927 -319 -907
rect -299 -927 -290 -907
rect -415 -935 -290 -927
rect -165 -965 -125 -950
rect -165 -985 -155 -965
rect -135 -985 -125 -965
rect 500 -959 535 -950
rect 560 -955 595 -900
rect 840 -875 880 -860
rect 840 -895 850 -875
rect 870 -895 880 -875
rect 840 -910 880 -895
rect 500 -976 512 -959
rect 529 -976 535 -959
rect 500 -985 535 -976
rect 550 -958 605 -955
rect 550 -975 569 -958
rect 586 -975 605 -958
rect 550 -980 605 -975
rect -165 -1000 -125 -985
rect 305 -1020 535 -985
rect 305 -1155 340 -1020
rect 830 -1030 880 -1020
rect 830 -1050 845 -1030
rect 865 -1050 880 -1030
rect 830 -1060 880 -1050
rect -70 -1190 340 -1155
rect -70 -1330 -35 -1190
rect 1020 -1315 1070 -1305
rect -70 -1337 75 -1330
rect -70 -1357 46 -1337
rect 66 -1357 75 -1337
rect 1020 -1335 1035 -1315
rect 1055 -1335 1070 -1315
rect 1020 -1345 1070 -1335
rect -70 -1370 75 -1357
rect -65 -1470 -25 -1455
rect -65 -1490 -55 -1470
rect -35 -1490 -25 -1470
rect -65 -1505 -25 -1490
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -348 0 1 -515
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1709947739
transform -1 0 1340 0 -1 -1281
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1709947739
transform 1 0 923 0 1 -1084
box -19 -24 203 296
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1709947739
transform 1 0 1140 0 1 -516
box -19 -24 203 296
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -7 0 1 -516
box -19 -24 985 296
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_1
timestamp 1709947739
transform -1 0 963 0 -1 -1281
box -19 -24 985 296
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 -336 0 1 -1037
box -19 -24 157 296
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1709947739
transform -1 0 -112 0 -1 -1281
box -19 -24 157 296
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 465 0 1 -1084
box -19 -24 341 296
<< end >>
