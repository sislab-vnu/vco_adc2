magic
tech sky130A
timestamp 1726647848
<< nwell >>
rect -130 -40 200 440
<< pmoshvt >>
rect 0 0 50 400
rect 90 0 140 400
<< pdiff >>
rect -40 390 0 400
rect -40 370 -30 390
rect -10 370 0 390
rect -40 350 0 370
rect -40 330 -30 350
rect -10 330 0 350
rect -40 310 0 330
rect -40 290 -30 310
rect -10 290 0 310
rect -40 270 0 290
rect -40 250 -30 270
rect -10 250 0 270
rect -40 230 0 250
rect -40 210 -30 230
rect -10 210 0 230
rect -40 190 0 210
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 390 90 400
rect 50 370 60 390
rect 80 370 90 390
rect 50 350 90 370
rect 50 330 60 350
rect 80 330 90 350
rect 50 310 90 330
rect 50 290 60 310
rect 80 290 90 310
rect 50 270 90 290
rect 50 250 60 270
rect 80 250 90 270
rect 50 230 90 250
rect 50 210 60 230
rect 80 210 90 230
rect 50 190 90 210
rect 50 170 60 190
rect 80 170 90 190
rect 50 150 90 170
rect 50 130 60 150
rect 80 130 90 150
rect 50 110 90 130
rect 50 90 60 110
rect 80 90 90 110
rect 50 70 90 90
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 390 180 400
rect 140 370 150 390
rect 170 370 180 390
rect 140 350 180 370
rect 140 330 150 350
rect 170 330 180 350
rect 140 310 180 330
rect 140 290 150 310
rect 170 290 180 310
rect 140 270 180 290
rect 140 250 150 270
rect 170 250 180 270
rect 140 230 180 250
rect 140 210 150 230
rect 170 210 180 230
rect 140 190 180 210
rect 140 170 150 190
rect 170 170 180 190
rect 140 150 180 170
rect 140 130 150 150
rect 170 130 180 150
rect 140 110 180 130
rect 140 90 150 110
rect 170 90 180 110
rect 140 70 180 90
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
<< pdiffc >>
rect -30 370 -10 390
rect -30 330 -10 350
rect -30 290 -10 310
rect -30 250 -10 270
rect -30 210 -10 230
rect -30 170 -10 190
rect -30 130 -10 150
rect -30 90 -10 110
rect -30 50 -10 70
rect -30 10 -10 30
rect 60 370 80 390
rect 60 330 80 350
rect 60 290 80 310
rect 60 250 80 270
rect 60 210 80 230
rect 60 170 80 190
rect 60 130 80 150
rect 60 90 80 110
rect 60 50 80 70
rect 60 10 80 30
rect 150 370 170 390
rect 150 330 170 350
rect 150 290 170 310
rect 150 250 170 270
rect 150 210 170 230
rect 150 170 170 190
rect 150 130 170 150
rect 150 90 170 110
rect 150 50 170 70
rect 150 10 170 30
<< nsubdiff >>
rect -110 390 -70 405
rect -110 370 -100 390
rect -80 370 -70 390
rect -110 355 -70 370
<< nsubdiffcont >>
rect -100 370 -80 390
<< poly >>
rect 0 475 140 490
rect 0 455 40 475
rect 100 455 140 475
rect 0 440 140 455
rect 0 400 50 440
rect 90 400 140 440
rect 0 -40 50 0
rect 90 -40 140 0
<< polycont >>
rect 40 455 100 475
<< locali >>
rect 25 475 115 490
rect 25 455 40 475
rect 100 455 115 475
rect 25 440 115 455
rect -110 390 -70 405
rect -110 370 -100 390
rect -80 370 -70 390
rect -110 355 -70 370
rect -40 390 0 400
rect -40 370 -30 390
rect -10 370 0 390
rect -40 350 0 370
rect -40 330 -30 350
rect -10 330 0 350
rect -40 310 0 330
rect -40 290 -30 310
rect -10 290 0 310
rect -40 270 0 290
rect -40 250 -30 270
rect -10 250 0 270
rect -40 230 0 250
rect -40 210 -30 230
rect -10 210 0 230
rect -40 190 0 210
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 390 90 400
rect 50 370 60 390
rect 80 370 90 390
rect 50 350 90 370
rect 50 330 60 350
rect 80 330 90 350
rect 50 310 90 330
rect 50 290 60 310
rect 80 290 90 310
rect 50 270 90 290
rect 50 250 60 270
rect 80 250 90 270
rect 50 230 90 250
rect 50 210 60 230
rect 80 210 90 230
rect 50 190 90 210
rect 50 170 60 190
rect 80 170 90 190
rect 50 150 90 170
rect 50 130 60 150
rect 80 130 90 150
rect 50 110 90 130
rect 50 90 60 110
rect 80 90 90 110
rect 50 70 90 90
rect 50 50 60 70
rect 80 50 90 70
rect 50 30 90 50
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
rect 140 390 180 400
rect 140 370 150 390
rect 170 370 180 390
rect 140 350 180 370
rect 140 330 150 350
rect 170 330 180 350
rect 140 310 180 330
rect 140 290 150 310
rect 170 290 180 310
rect 140 270 180 290
rect 140 250 150 270
rect 170 250 180 270
rect 140 230 180 250
rect 140 210 150 230
rect 170 210 180 230
rect 140 190 180 210
rect 140 170 150 190
rect 170 170 180 190
rect 140 150 180 170
rect 140 130 150 150
rect 170 130 180 150
rect 140 110 180 130
rect 140 90 150 110
rect 170 90 180 110
rect 140 70 180 90
rect 140 50 150 70
rect 170 50 180 70
rect 140 30 180 50
rect 140 10 150 30
rect 170 10 180 30
rect 140 0 180 10
<< viali >>
rect 40 455 100 475
rect -100 370 -80 390
rect -30 370 -10 390
rect -30 330 -10 350
rect -30 50 -10 70
rect -30 10 -10 30
rect 150 370 170 390
rect 150 330 170 350
rect 150 50 170 70
rect 150 10 170 30
<< metal1 >>
rect 0 475 140 490
rect 0 455 40 475
rect 100 455 140 475
rect 0 440 140 455
rect -110 390 -70 405
rect -110 370 -100 390
rect -80 370 -70 390
rect -110 355 -70 370
rect -40 390 0 400
rect -40 370 -30 390
rect -10 385 0 390
rect 140 390 180 400
rect 140 385 150 390
rect -10 370 150 385
rect 170 370 180 390
rect -40 350 180 370
rect -40 330 -30 350
rect -10 335 150 350
rect -10 330 0 335
rect -40 320 0 330
rect 140 330 150 335
rect 170 330 180 350
rect 140 320 180 330
rect -40 70 0 80
rect -40 50 -30 70
rect -10 65 0 70
rect 140 70 180 80
rect 140 65 150 70
rect -10 50 150 65
rect 170 50 180 70
rect -40 30 180 50
rect -40 10 -30 30
rect -10 15 150 30
rect -10 10 0 15
rect -40 0 0 10
rect 140 10 150 15
rect 170 10 180 30
rect 140 0 180 10
<< labels >>
rlabel metal1 -90 405 -90 405 1 B
port 4 n
rlabel metal1 -20 400 -20 400 1 S
port 2 n
rlabel locali 70 0 70 0 5 D
port 3 s
rlabel metal1 70 490 70 490 1 G
port 1 n
<< end >>
