* NGSPICE file created from x5s_cc_osc.ext - technology: sky130A

.subckt aux_inv A Y VGND VDDA GND
X0 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=2 ps=10.8 w=5 l=3.65
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=1.6 ps=8.8 w=4 l=3.65
.ends

.subckt main_inv A Y VGND GND VDDA
X0 VDDA A Y VDDA sky130_fd_pr__pfet_01v8 ad=2 pd=10.8 as=1 ps=5.4 w=5 l=3.65 M=2
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=3.65 M=2
.ends

.subckt cc_inv inp inn outp outn VGND GND VDDA
Xaux_inv_0 outp outn VGND VDDA GND aux_inv
Xaux_inv_1 outn outp VGND VDDA GND aux_inv
Xmain_inv_0 inp outp VGND GND VDDA main_inv
Xmain_inv_1 inn outn VGND GND VDDA main_inv
.ends

.subckt x5s_cc_osc pn[0] pn[1] pn[2] pn[3] pn[4] p[0] p[1] p[2] p[3] p[4] VGND VDDA
+ GND
Xcc_inv_0 p[4] pn[4] p[0] pn[0] VGND GND VDDA cc_inv
Xcc_inv_2 p[1] pn[1] p[2] pn[2] VGND GND VDDA cc_inv
Xcc_inv_1 p[0] pn[0] p[1] pn[1] VGND GND VDDA cc_inv
Xcc_inv_3 p[3] pn[3] p[4] pn[4] VGND GND VDDA cc_inv
Xcc_inv_4 p[2] pn[2] p[3] pn[3] VGND GND VDDA cc_inv
.ends


