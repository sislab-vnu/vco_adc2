magic
tech sky130A
timestamp 1724146945
<< pwell >>
rect -60 -40 830 440
<< nmos >>
rect 0 0 365 400
rect 405 0 770 400
<< ndiff >>
rect -40 390 0 400
rect -40 370 -30 390
rect -10 370 0 390
rect -40 350 0 370
rect -40 330 -30 350
rect -10 330 0 350
rect -40 310 0 330
rect -40 290 -30 310
rect -10 290 0 310
rect -40 270 0 290
rect -40 250 -30 270
rect -10 250 0 270
rect -40 230 0 250
rect -40 210 -30 230
rect -10 210 0 230
rect -40 190 0 210
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 365 390 405 400
rect 365 370 375 390
rect 395 370 405 390
rect 365 350 405 370
rect 365 330 375 350
rect 395 330 405 350
rect 365 310 405 330
rect 365 290 375 310
rect 395 290 405 310
rect 365 270 405 290
rect 365 250 375 270
rect 395 250 405 270
rect 365 230 405 250
rect 365 210 375 230
rect 395 210 405 230
rect 365 190 405 210
rect 365 170 375 190
rect 395 170 405 190
rect 365 150 405 170
rect 365 130 375 150
rect 395 130 405 150
rect 365 110 405 130
rect 365 90 375 110
rect 395 90 405 110
rect 365 70 405 90
rect 365 50 375 70
rect 395 50 405 70
rect 365 30 405 50
rect 365 10 375 30
rect 395 10 405 30
rect 365 0 405 10
rect 770 390 810 400
rect 770 370 780 390
rect 800 370 810 390
rect 770 350 810 370
rect 770 330 780 350
rect 800 330 810 350
rect 770 310 810 330
rect 770 290 780 310
rect 800 290 810 310
rect 770 270 810 290
rect 770 250 780 270
rect 800 250 810 270
rect 770 230 810 250
rect 770 210 780 230
rect 800 210 810 230
rect 770 190 810 210
rect 770 170 780 190
rect 800 170 810 190
rect 770 150 810 170
rect 770 130 780 150
rect 800 130 810 150
rect 770 110 810 130
rect 770 90 780 110
rect 800 90 810 110
rect 770 70 810 90
rect 770 50 780 70
rect 800 50 810 70
rect 770 30 810 50
rect 770 10 780 30
rect 800 10 810 30
rect 770 0 810 10
<< ndiffc >>
rect -30 370 -10 390
rect -30 330 -10 350
rect -30 290 -10 310
rect -30 250 -10 270
rect -30 210 -10 230
rect -30 170 -10 190
rect -30 130 -10 150
rect -30 90 -10 110
rect -30 50 -10 70
rect -30 10 -10 30
rect 375 370 395 390
rect 375 330 395 350
rect 375 290 395 310
rect 375 250 395 270
rect 375 210 395 230
rect 375 170 395 190
rect 375 130 395 150
rect 375 90 395 110
rect 375 50 395 70
rect 375 10 395 30
rect 780 370 800 390
rect 780 330 800 350
rect 780 290 800 310
rect 780 250 800 270
rect 780 210 800 230
rect 780 170 800 190
rect 780 130 800 150
rect 780 90 800 110
rect 780 50 800 70
rect 780 10 800 30
<< poly >>
rect 0 400 365 440
rect 405 400 770 440
rect 0 -40 365 0
rect 405 -40 770 0
<< locali >>
rect -40 390 0 400
rect -40 370 -30 390
rect -10 370 0 390
rect -40 350 0 370
rect -40 330 -30 350
rect -10 330 0 350
rect -40 310 0 330
rect -40 290 -30 310
rect -10 290 0 310
rect -40 270 0 290
rect -40 250 -30 270
rect -10 250 0 270
rect -40 230 0 250
rect -40 210 -30 230
rect -10 210 0 230
rect -40 190 0 210
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 365 390 405 400
rect 365 370 375 390
rect 395 370 405 390
rect 365 350 405 370
rect 365 330 375 350
rect 395 330 405 350
rect 365 310 405 330
rect 365 290 375 310
rect 395 290 405 310
rect 365 270 405 290
rect 365 250 375 270
rect 395 250 405 270
rect 365 230 405 250
rect 365 210 375 230
rect 395 210 405 230
rect 365 190 405 210
rect 365 170 375 190
rect 395 170 405 190
rect 365 150 405 170
rect 365 130 375 150
rect 395 130 405 150
rect 365 110 405 130
rect 365 90 375 110
rect 395 90 405 110
rect 365 70 405 90
rect 365 50 375 70
rect 395 50 405 70
rect 365 30 405 50
rect 365 10 375 30
rect 395 10 405 30
rect 365 0 405 10
rect 770 390 810 400
rect 770 370 780 390
rect 800 370 810 390
rect 770 350 810 370
rect 770 330 780 350
rect 800 330 810 350
rect 770 310 810 330
rect 770 290 780 310
rect 800 290 810 310
rect 770 270 810 290
rect 770 250 780 270
rect 800 250 810 270
rect 770 230 810 250
rect 770 210 780 230
rect 800 210 810 230
rect 770 190 810 210
rect 770 170 780 190
rect 800 170 810 190
rect 770 150 810 170
rect 770 130 780 150
rect 800 130 810 150
rect 770 110 810 130
rect 770 90 780 110
rect 800 90 810 110
rect 770 70 810 90
rect 770 50 780 70
rect 800 50 810 70
rect 770 30 810 50
rect 770 10 780 30
rect 800 10 810 30
rect 770 0 810 10
<< labels >>
rlabel locali -20 400 -20 400 1 S
port 1 n
rlabel locali 385 400 385 400 1 D
port 2 n
rlabel locali 790 400 790 400 1 S
port 3 n
rlabel poly 170 -40 170 -40 5 G
port 4 s
rlabel poly 590 -40 590 -40 5 G
port 5 s
<< end >>
